.SUBCKT layer1 vdd vss in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15 in16 in17 in18 in19 in20 in21 in22 in23 in24 in25 in26 in27 in28 in29 in30 in31 in32 in33 in34 in35 in36 in37 in38 in39 in40 in41 in42 in43 in44 in45 in46 in47 in48 in49 in50 in51 in52 in53 in54 in55 in56 in57 in58 in59 in60 in61 in62 in63 in64 in65 in66 in67 in68 in69 in70 in71 in72 in73 in74 in75 in76 in77 in78 in79 in80 in81 in82 in83 in84 in85 in86 in87 in88 in89 in90 in91 in92 in93 in94 in95 in96 in97 in98 in99 in100 in101 in102 in103 in104 in105 in106 in107 in108 in109 in110 in111 in112 in113 in114 in115 in116 in117 in118 in119 in120 in121 in122 in123 in124 in125 in126 in127 in128 in129 in130 in131 in132 in133 in134 in135 in136 in137 in138 in139 in140 in141 in142 in143 in144 in145 in146 in147 in148 in149 in150 in151 in152 in153 in154 in155 in156 in157 in158 in159 in160 in161 in162 in163 in164 in165 in166 in167 in168 in169 in170 in171 in172 in173 in174 in175 in176 in177 in178 in179 in180 in181 in182 in183 in184 in185 in186 in187 in188 in189 in190 in191 in192 in193 in194 in195 in196 in197 in198 in199 in200 in201 in202 in203 in204 in205 in206 in207 in208 in209 in210 in211 in212 in213 in214 in215 in216 in217 in218 in219 in220 in221 in222 in223 in224 in225 in226 in227 in228 in229 in230 in231 in232 in233 in234 in235 in236 in237 in238 in239 in240 in241 in242 in243 in244 in245 in246 in247 in248 in249 in250 in251 in252 in253 in254 in255 in256 in257 in258 in259 in260 in261 in262 in263 in264 in265 in266 in267 in268 in269 in270 in271 in272 in273 in274 in275 in276 in277 in278 in279 in280 in281 in282 in283 in284 in285 in286 in287 in288 in289 in290 in291 in292 in293 in294 in295 in296 in297 in298 in299 in300 in301 in302 in303 in304 in305 in306 in307 in308 in309 in310 in311 in312 in313 in314 in315 in316 in317 in318 in319 in320 in321 in322 in323 in324 in325 in326 in327 in328 in329 in330 in331 in332 in333 in334 in335 in336 in337 in338 in339 in340 in341 in342 in343 in344 in345 in346 in347 in348 in349 in350 in351 in352 in353 in354 in355 in356 in357 in358 in359 in360 in361 in362 in363 in364 in365 in366 in367 in368 in369 in370 in371 in372 in373 in374 in375 in376 in377 in378 in379 in380 in381 in382 in383 in384 in385 in386 in387 in388 in389 in390 in391 in392 in393 in394 in395 in396 in397 in398 in399 in400 in401 in402 in403 in404 in405 in406 in407 in408 in409 in410 in411 in412 in413 in414 in415 in416 in417 in418 in419 in420 in421 in422 in423 in424 in425 in426 in427 in428 in429 in430 in431 in432 in433 in434 in435 in436 in437 in438 in439 in440 in441 in442 in443 in444 in445 in446 in447 in448 in449 in450 in451 in452 in453 in454 in455 in456 in457 in458 in459 in460 in461 in462 in463 in464 in465 in466 in467 in468 in469 in470 in471 in472 in473 in474 in475 in476 in477 in478 in479 in480 in481 in482 in483 in484 in485 in486 in487 in488 in489 in490 in491 in492 in493 in494 in495 in496 in497 in498 in499 in500 in501 in502 in503 in504 in505 in506 in507 in508 in509 in510 in511 in512 in513 in514 in515 in516 in517 in518 in519 in520 in521 in522 in523 in524 in525 in526 in527 in528 in529 in530 in531 in532 in533 in534 in535 in536 in537 in538 in539 in540 in541 in542 in543 in544 in545 in546 in547 in548 in549 in550 in551 in552 in553 in554 in555 in556 in557 in558 in559 in560 in561 in562 in563 in564 in565 in566 in567 in568 in569 in570 in571 in572 in573 in574 in575 in576 in577 in578 in579 in580 in581 in582 in583 in584 in585 in586 in587 in588 in589 in590 in591 in592 in593 in594 in595 in596 in597 in598 in599 in600 in601 in602 in603 in604 in605 in606 in607 in608 in609 in610 in611 in612 in613 in614 in615 in616 in617 in618 in619 in620 in621 in622 in623 in624 in625 in626 in627 in628 in629 in630 in631 in632 in633 in634 in635 in636 in637 in638 in639 in640 in641 in642 in643 in644 in645 in646 in647 in648 in649 in650 in651 in652 in653 in654 in655 in656 in657 in658 in659 in660 in661 in662 in663 in664 in665 in666 in667 in668 in669 in670 in671 in672 in673 in674 in675 in676 in677 in678 in679 in680 in681 in682 in683 in684 in685 in686 in687 in688 in689 in690 in691 in692 in693 in694 in695 in696 in697 in698 in699 in700 in701 in702 in703 in704 in705 in706 in707 in708 in709 in710 in711 in712 in713 in714 in715 in716 in717 in718 in719 in720 in721 in722 in723 in724 in725 in726 in727 in728 in729 in730 in731 in732 in733 in734 in735 in736 in737 in738 in739 in740 in741 in742 in743 in744 in745 in746 in747 in748 in749 in750 in751 in752 in753 in754 in755 in756 in757 in758 in759 in760 in761 in762 in763 in764 in765 in766 in767 in768 in769 in770 in771 in772 in773 in774 in775 in776 in777 in778 in779 in780 in781 in782 in783 in784 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 out11 out12 out13 out14 out15 out16 out17 out18 out19 out20 out21 out22 out23 out24 out25 out26 out27 out28 out29 out30 out31 out32 out33 out34 out35 out36 out37 out38 out39 out40 out41 out42 out43 out44 out45 out46 out47 out48 out49 out50 out51 out52 out53 out54 out55 out56 out57 out58 out59 out60 out61 out62 out63 out64 out65 out66 out67 out68 out69 out70 out71 out72 out73 out74 out75 out76 out77 out78 out79 out80 out81 out82 out83 out84 out85 out86 out87 out88 out89 out90 out91 out92 out93 out94 out95 out96 out97 out98 out99 out100 

**********Non-Negative Weighted Array****************
Rwpos1_1 in1 sp1 11140.846016
Rwpos1_2 in1 sp2 3183.098862
Rwpos1_3 in1 sp3 3183.098862
Rwpos1_4 in1 sp4 3183.098862
Rwpos1_5 in1 sp5 11140.846016
Rwpos1_6 in1 sp6 3183.098862
Rwpos1_7 in1 sp7 3183.098862
Rwpos1_8 in1 sp8 11140.846016
Rwpos1_9 in1 sp9 11140.846016
Rwpos1_10 in1 sp10 3183.098862
Rwpos1_11 in1 sp11 11140.846016
Rwpos1_12 in1 sp12 3183.098862
Rwpos1_13 in1 sp13 3183.098862
Rwpos1_14 in1 sp14 3183.098862
Rwpos1_15 in1 sp15 11140.846016
Rwpos1_16 in1 sp16 3183.098862
Rwpos1_17 in1 sp17 11140.846016
Rwpos1_18 in1 sp18 11140.846016
Rwpos1_19 in1 sp19 3183.098862
Rwpos1_20 in1 sp20 3183.098862
Rwpos1_21 in1 sp21 3183.098862
Rwpos1_22 in1 sp22 3183.098862
Rwpos1_23 in1 sp23 3183.098862
Rwpos1_24 in1 sp24 3183.098862
Rwpos1_25 in1 sp25 11140.846016
Rwpos1_26 in1 sp26 3183.098862
Rwpos1_27 in1 sp27 3183.098862
Rwpos1_28 in1 sp28 11140.846016
Rwpos1_29 in1 sp29 11140.846016
Rwpos1_30 in1 sp30 3183.098862
Rwpos1_31 in1 sp31 11140.846016
Rwpos1_32 in1 sp32 3183.098862
Rwpos1_33 in1 sp33 11140.846016
Rwpos1_34 in1 sp34 3183.098862
Rwpos1_35 in1 sp35 3183.098862
Rwpos1_36 in1 sp36 11140.846016
Rwpos1_37 in1 sp37 3183.098862
Rwpos1_38 in1 sp38 3183.098862
Rwpos1_39 in1 sp39 11140.846016
Rwpos1_40 in1 sp40 11140.846016
Rwpos1_41 in1 sp41 3183.098862
Rwpos1_42 in1 sp42 3183.098862
Rwpos1_43 in1 sp43 3183.098862
Rwpos1_44 in1 sp44 11140.846016
Rwpos1_45 in1 sp45 11140.846016
Rwpos1_46 in1 sp46 3183.098862
Rwpos1_47 in1 sp47 11140.846016
Rwpos1_48 in1 sp48 11140.846016
Rwpos1_49 in1 sp49 3183.098862
Rwpos1_50 in1 sp50 3183.098862
Rwpos1_51 in1 sp51 3183.098862
Rwpos1_52 in1 sp52 11140.846016
Rwpos1_53 in1 sp53 11140.846016
Rwpos1_54 in1 sp54 11140.846016
Rwpos1_55 in1 sp55 3183.098862
Rwpos1_56 in1 sp56 3183.098862
Rwpos1_57 in1 sp57 11140.846016
Rwpos1_58 in1 sp58 3183.098862
Rwpos1_59 in1 sp59 11140.846016
Rwpos1_60 in1 sp60 3183.098862
Rwpos1_61 in1 sp61 3183.098862
Rwpos1_62 in1 sp62 11140.846016
Rwpos1_63 in1 sp63 3183.098862
Rwpos1_64 in1 sp64 3183.098862
Rwpos1_65 in1 sp65 11140.846016
Rwpos1_66 in1 sp66 11140.846016
Rwpos1_67 in1 sp67 3183.098862
Rwpos1_68 in1 sp68 11140.846016
Rwpos1_69 in1 sp69 11140.846016
Rwpos1_70 in1 sp70 3183.098862
Rwpos1_71 in1 sp71 11140.846016
Rwpos1_72 in1 sp72 11140.846016
Rwpos1_73 in1 sp73 11140.846016
Rwpos1_74 in1 sp74 3183.098862
Rwpos1_75 in1 sp75 3183.098862
Rwpos1_76 in1 sp76 3183.098862
Rwpos1_77 in1 sp77 3183.098862
Rwpos1_78 in1 sp78 11140.846016
Rwpos1_79 in1 sp79 11140.846016
Rwpos1_80 in1 sp80 11140.846016
Rwpos1_81 in1 sp81 11140.846016
Rwpos1_82 in1 sp82 3183.098862
Rwpos1_83 in1 sp83 11140.846016
Rwpos1_84 in1 sp84 11140.846016
Rwpos1_85 in1 sp85 11140.846016
Rwpos1_86 in1 sp86 11140.846016
Rwpos1_87 in1 sp87 11140.846016
Rwpos1_88 in1 sp88 11140.846016
Rwpos1_89 in1 sp89 11140.846016
Rwpos1_90 in1 sp90 11140.846016
Rwpos1_91 in1 sp91 11140.846016
Rwpos1_92 in1 sp92 3183.098862
Rwpos1_93 in1 sp93 3183.098862
Rwpos1_94 in1 sp94 11140.846016
Rwpos1_95 in1 sp95 3183.098862
Rwpos1_96 in1 sp96 11140.846016
Rwpos1_97 in1 sp97 11140.846016
Rwpos1_98 in1 sp98 11140.846016
Rwpos1_99 in1 sp99 3183.098862
Rwpos1_100 in1 sp100 3183.098862
Rwpos2_1 in2 sp1 3183.098862
Rwpos2_2 in2 sp2 3183.098862
Rwpos2_3 in2 sp3 11140.846016
Rwpos2_4 in2 sp4 3183.098862
Rwpos2_5 in2 sp5 3183.098862
Rwpos2_6 in2 sp6 11140.846016
Rwpos2_7 in2 sp7 11140.846016
Rwpos2_8 in2 sp8 3183.098862
Rwpos2_9 in2 sp9 11140.846016
Rwpos2_10 in2 sp10 3183.098862
Rwpos2_11 in2 sp11 3183.098862
Rwpos2_12 in2 sp12 3183.098862
Rwpos2_13 in2 sp13 11140.846016
Rwpos2_14 in2 sp14 3183.098862
Rwpos2_15 in2 sp15 11140.846016
Rwpos2_16 in2 sp16 11140.846016
Rwpos2_17 in2 sp17 3183.098862
Rwpos2_18 in2 sp18 3183.098862
Rwpos2_19 in2 sp19 11140.846016
Rwpos2_20 in2 sp20 11140.846016
Rwpos2_21 in2 sp21 3183.098862
Rwpos2_22 in2 sp22 3183.098862
Rwpos2_23 in2 sp23 11140.846016
Rwpos2_24 in2 sp24 11140.846016
Rwpos2_25 in2 sp25 3183.098862
Rwpos2_26 in2 sp26 11140.846016
Rwpos2_27 in2 sp27 3183.098862
Rwpos2_28 in2 sp28 3183.098862
Rwpos2_29 in2 sp29 11140.846016
Rwpos2_30 in2 sp30 3183.098862
Rwpos2_31 in2 sp31 3183.098862
Rwpos2_32 in2 sp32 3183.098862
Rwpos2_33 in2 sp33 3183.098862
Rwpos2_34 in2 sp34 3183.098862
Rwpos2_35 in2 sp35 3183.098862
Rwpos2_36 in2 sp36 11140.846016
Rwpos2_37 in2 sp37 11140.846016
Rwpos2_38 in2 sp38 11140.846016
Rwpos2_39 in2 sp39 3183.098862
Rwpos2_40 in2 sp40 3183.098862
Rwpos2_41 in2 sp41 11140.846016
Rwpos2_42 in2 sp42 11140.846016
Rwpos2_43 in2 sp43 3183.098862
Rwpos2_44 in2 sp44 11140.846016
Rwpos2_45 in2 sp45 11140.846016
Rwpos2_46 in2 sp46 3183.098862
Rwpos2_47 in2 sp47 11140.846016
Rwpos2_48 in2 sp48 11140.846016
Rwpos2_49 in2 sp49 3183.098862
Rwpos2_50 in2 sp50 11140.846016
Rwpos2_51 in2 sp51 3183.098862
Rwpos2_52 in2 sp52 11140.846016
Rwpos2_53 in2 sp53 11140.846016
Rwpos2_54 in2 sp54 3183.098862
Rwpos2_55 in2 sp55 3183.098862
Rwpos2_56 in2 sp56 11140.846016
Rwpos2_57 in2 sp57 11140.846016
Rwpos2_58 in2 sp58 3183.098862
Rwpos2_59 in2 sp59 11140.846016
Rwpos2_60 in2 sp60 11140.846016
Rwpos2_61 in2 sp61 11140.846016
Rwpos2_62 in2 sp62 11140.846016
Rwpos2_63 in2 sp63 11140.846016
Rwpos2_64 in2 sp64 11140.846016
Rwpos2_65 in2 sp65 3183.098862
Rwpos2_66 in2 sp66 11140.846016
Rwpos2_67 in2 sp67 11140.846016
Rwpos2_68 in2 sp68 11140.846016
Rwpos2_69 in2 sp69 11140.846016
Rwpos2_70 in2 sp70 11140.846016
Rwpos2_71 in2 sp71 3183.098862
Rwpos2_72 in2 sp72 11140.846016
Rwpos2_73 in2 sp73 11140.846016
Rwpos2_74 in2 sp74 11140.846016
Rwpos2_75 in2 sp75 11140.846016
Rwpos2_76 in2 sp76 11140.846016
Rwpos2_77 in2 sp77 3183.098862
Rwpos2_78 in2 sp78 3183.098862
Rwpos2_79 in2 sp79 11140.846016
Rwpos2_80 in2 sp80 3183.098862
Rwpos2_81 in2 sp81 3183.098862
Rwpos2_82 in2 sp82 11140.846016
Rwpos2_83 in2 sp83 11140.846016
Rwpos2_84 in2 sp84 3183.098862
Rwpos2_85 in2 sp85 3183.098862
Rwpos2_86 in2 sp86 11140.846016
Rwpos2_87 in2 sp87 11140.846016
Rwpos2_88 in2 sp88 11140.846016
Rwpos2_89 in2 sp89 3183.098862
Rwpos2_90 in2 sp90 11140.846016
Rwpos2_91 in2 sp91 3183.098862
Rwpos2_92 in2 sp92 3183.098862
Rwpos2_93 in2 sp93 3183.098862
Rwpos2_94 in2 sp94 3183.098862
Rwpos2_95 in2 sp95 11140.846016
Rwpos2_96 in2 sp96 3183.098862
Rwpos2_97 in2 sp97 11140.846016
Rwpos2_98 in2 sp98 11140.846016
Rwpos2_99 in2 sp99 11140.846016
Rwpos2_100 in2 sp100 11140.846016
Rwpos3_1 in3 sp1 3183.098862
Rwpos3_2 in3 sp2 11140.846016
Rwpos3_3 in3 sp3 11140.846016
Rwpos3_4 in3 sp4 3183.098862
Rwpos3_5 in3 sp5 11140.846016
Rwpos3_6 in3 sp6 11140.846016
Rwpos3_7 in3 sp7 3183.098862
Rwpos3_8 in3 sp8 11140.846016
Rwpos3_9 in3 sp9 11140.846016
Rwpos3_10 in3 sp10 11140.846016
Rwpos3_11 in3 sp11 11140.846016
Rwpos3_12 in3 sp12 3183.098862
Rwpos3_13 in3 sp13 3183.098862
Rwpos3_14 in3 sp14 11140.846016
Rwpos3_15 in3 sp15 3183.098862
Rwpos3_16 in3 sp16 3183.098862
Rwpos3_17 in3 sp17 3183.098862
Rwpos3_18 in3 sp18 3183.098862
Rwpos3_19 in3 sp19 3183.098862
Rwpos3_20 in3 sp20 11140.846016
Rwpos3_21 in3 sp21 3183.098862
Rwpos3_22 in3 sp22 3183.098862
Rwpos3_23 in3 sp23 3183.098862
Rwpos3_24 in3 sp24 11140.846016
Rwpos3_25 in3 sp25 11140.846016
Rwpos3_26 in3 sp26 11140.846016
Rwpos3_27 in3 sp27 11140.846016
Rwpos3_28 in3 sp28 11140.846016
Rwpos3_29 in3 sp29 11140.846016
Rwpos3_30 in3 sp30 3183.098862
Rwpos3_31 in3 sp31 11140.846016
Rwpos3_32 in3 sp32 3183.098862
Rwpos3_33 in3 sp33 3183.098862
Rwpos3_34 in3 sp34 3183.098862
Rwpos3_35 in3 sp35 11140.846016
Rwpos3_36 in3 sp36 3183.098862
Rwpos3_37 in3 sp37 11140.846016
Rwpos3_38 in3 sp38 11140.846016
Rwpos3_39 in3 sp39 11140.846016
Rwpos3_40 in3 sp40 3183.098862
Rwpos3_41 in3 sp41 11140.846016
Rwpos3_42 in3 sp42 11140.846016
Rwpos3_43 in3 sp43 3183.098862
Rwpos3_44 in3 sp44 11140.846016
Rwpos3_45 in3 sp45 3183.098862
Rwpos3_46 in3 sp46 11140.846016
Rwpos3_47 in3 sp47 3183.098862
Rwpos3_48 in3 sp48 11140.846016
Rwpos3_49 in3 sp49 3183.098862
Rwpos3_50 in3 sp50 11140.846016
Rwpos3_51 in3 sp51 3183.098862
Rwpos3_52 in3 sp52 11140.846016
Rwpos3_53 in3 sp53 3183.098862
Rwpos3_54 in3 sp54 3183.098862
Rwpos3_55 in3 sp55 11140.846016
Rwpos3_56 in3 sp56 11140.846016
Rwpos3_57 in3 sp57 3183.098862
Rwpos3_58 in3 sp58 11140.846016
Rwpos3_59 in3 sp59 3183.098862
Rwpos3_60 in3 sp60 11140.846016
Rwpos3_61 in3 sp61 3183.098862
Rwpos3_62 in3 sp62 11140.846016
Rwpos3_63 in3 sp63 3183.098862
Rwpos3_64 in3 sp64 11140.846016
Rwpos3_65 in3 sp65 3183.098862
Rwpos3_66 in3 sp66 3183.098862
Rwpos3_67 in3 sp67 3183.098862
Rwpos3_68 in3 sp68 11140.846016
Rwpos3_69 in3 sp69 3183.098862
Rwpos3_70 in3 sp70 3183.098862
Rwpos3_71 in3 sp71 3183.098862
Rwpos3_72 in3 sp72 11140.846016
Rwpos3_73 in3 sp73 3183.098862
Rwpos3_74 in3 sp74 11140.846016
Rwpos3_75 in3 sp75 3183.098862
Rwpos3_76 in3 sp76 11140.846016
Rwpos3_77 in3 sp77 11140.846016
Rwpos3_78 in3 sp78 3183.098862
Rwpos3_79 in3 sp79 11140.846016
Rwpos3_80 in3 sp80 11140.846016
Rwpos3_81 in3 sp81 11140.846016
Rwpos3_82 in3 sp82 3183.098862
Rwpos3_83 in3 sp83 3183.098862
Rwpos3_84 in3 sp84 11140.846016
Rwpos3_85 in3 sp85 3183.098862
Rwpos3_86 in3 sp86 3183.098862
Rwpos3_87 in3 sp87 11140.846016
Rwpos3_88 in3 sp88 3183.098862
Rwpos3_89 in3 sp89 11140.846016
Rwpos3_90 in3 sp90 3183.098862
Rwpos3_91 in3 sp91 3183.098862
Rwpos3_92 in3 sp92 3183.098862
Rwpos3_93 in3 sp93 11140.846016
Rwpos3_94 in3 sp94 11140.846016
Rwpos3_95 in3 sp95 3183.098862
Rwpos3_96 in3 sp96 11140.846016
Rwpos3_97 in3 sp97 11140.846016
Rwpos3_98 in3 sp98 3183.098862
Rwpos3_99 in3 sp99 3183.098862
Rwpos3_100 in3 sp100 11140.846016
Rwpos4_1 in4 sp1 3183.098862
Rwpos4_2 in4 sp2 3183.098862
Rwpos4_3 in4 sp3 11140.846016
Rwpos4_4 in4 sp4 3183.098862
Rwpos4_5 in4 sp5 3183.098862
Rwpos4_6 in4 sp6 11140.846016
Rwpos4_7 in4 sp7 11140.846016
Rwpos4_8 in4 sp8 3183.098862
Rwpos4_9 in4 sp9 11140.846016
Rwpos4_10 in4 sp10 11140.846016
Rwpos4_11 in4 sp11 3183.098862
Rwpos4_12 in4 sp12 11140.846016
Rwpos4_13 in4 sp13 11140.846016
Rwpos4_14 in4 sp14 11140.846016
Rwpos4_15 in4 sp15 3183.098862
Rwpos4_16 in4 sp16 11140.846016
Rwpos4_17 in4 sp17 3183.098862
Rwpos4_18 in4 sp18 11140.846016
Rwpos4_19 in4 sp19 3183.098862
Rwpos4_20 in4 sp20 11140.846016
Rwpos4_21 in4 sp21 11140.846016
Rwpos4_22 in4 sp22 11140.846016
Rwpos4_23 in4 sp23 11140.846016
Rwpos4_24 in4 sp24 3183.098862
Rwpos4_25 in4 sp25 11140.846016
Rwpos4_26 in4 sp26 3183.098862
Rwpos4_27 in4 sp27 3183.098862
Rwpos4_28 in4 sp28 3183.098862
Rwpos4_29 in4 sp29 11140.846016
Rwpos4_30 in4 sp30 11140.846016
Rwpos4_31 in4 sp31 3183.098862
Rwpos4_32 in4 sp32 11140.846016
Rwpos4_33 in4 sp33 3183.098862
Rwpos4_34 in4 sp34 3183.098862
Rwpos4_35 in4 sp35 11140.846016
Rwpos4_36 in4 sp36 3183.098862
Rwpos4_37 in4 sp37 3183.098862
Rwpos4_38 in4 sp38 3183.098862
Rwpos4_39 in4 sp39 3183.098862
Rwpos4_40 in4 sp40 11140.846016
Rwpos4_41 in4 sp41 11140.846016
Rwpos4_42 in4 sp42 11140.846016
Rwpos4_43 in4 sp43 3183.098862
Rwpos4_44 in4 sp44 11140.846016
Rwpos4_45 in4 sp45 11140.846016
Rwpos4_46 in4 sp46 11140.846016
Rwpos4_47 in4 sp47 3183.098862
Rwpos4_48 in4 sp48 11140.846016
Rwpos4_49 in4 sp49 3183.098862
Rwpos4_50 in4 sp50 3183.098862
Rwpos4_51 in4 sp51 3183.098862
Rwpos4_52 in4 sp52 3183.098862
Rwpos4_53 in4 sp53 3183.098862
Rwpos4_54 in4 sp54 3183.098862
Rwpos4_55 in4 sp55 11140.846016
Rwpos4_56 in4 sp56 11140.846016
Rwpos4_57 in4 sp57 11140.846016
Rwpos4_58 in4 sp58 3183.098862
Rwpos4_59 in4 sp59 11140.846016
Rwpos4_60 in4 sp60 11140.846016
Rwpos4_61 in4 sp61 3183.098862
Rwpos4_62 in4 sp62 11140.846016
Rwpos4_63 in4 sp63 11140.846016
Rwpos4_64 in4 sp64 3183.098862
Rwpos4_65 in4 sp65 3183.098862
Rwpos4_66 in4 sp66 11140.846016
Rwpos4_67 in4 sp67 11140.846016
Rwpos4_68 in4 sp68 3183.098862
Rwpos4_69 in4 sp69 3183.098862
Rwpos4_70 in4 sp70 3183.098862
Rwpos4_71 in4 sp71 11140.846016
Rwpos4_72 in4 sp72 3183.098862
Rwpos4_73 in4 sp73 3183.098862
Rwpos4_74 in4 sp74 11140.846016
Rwpos4_75 in4 sp75 11140.846016
Rwpos4_76 in4 sp76 3183.098862
Rwpos4_77 in4 sp77 11140.846016
Rwpos4_78 in4 sp78 3183.098862
Rwpos4_79 in4 sp79 11140.846016
Rwpos4_80 in4 sp80 3183.098862
Rwpos4_81 in4 sp81 3183.098862
Rwpos4_82 in4 sp82 3183.098862
Rwpos4_83 in4 sp83 11140.846016
Rwpos4_84 in4 sp84 11140.846016
Rwpos4_85 in4 sp85 11140.846016
Rwpos4_86 in4 sp86 11140.846016
Rwpos4_87 in4 sp87 3183.098862
Rwpos4_88 in4 sp88 3183.098862
Rwpos4_89 in4 sp89 3183.098862
Rwpos4_90 in4 sp90 3183.098862
Rwpos4_91 in4 sp91 3183.098862
Rwpos4_92 in4 sp92 3183.098862
Rwpos4_93 in4 sp93 11140.846016
Rwpos4_94 in4 sp94 3183.098862
Rwpos4_95 in4 sp95 3183.098862
Rwpos4_96 in4 sp96 3183.098862
Rwpos4_97 in4 sp97 11140.846016
Rwpos4_98 in4 sp98 11140.846016
Rwpos4_99 in4 sp99 3183.098862
Rwpos4_100 in4 sp100 11140.846016
Rwpos5_1 in5 sp1 11140.846016
Rwpos5_2 in5 sp2 11140.846016
Rwpos5_3 in5 sp3 3183.098862
Rwpos5_4 in5 sp4 11140.846016
Rwpos5_5 in5 sp5 3183.098862
Rwpos5_6 in5 sp6 3183.098862
Rwpos5_7 in5 sp7 11140.846016
Rwpos5_8 in5 sp8 11140.846016
Rwpos5_9 in5 sp9 3183.098862
Rwpos5_10 in5 sp10 11140.846016
Rwpos5_11 in5 sp11 11140.846016
Rwpos5_12 in5 sp12 3183.098862
Rwpos5_13 in5 sp13 3183.098862
Rwpos5_14 in5 sp14 3183.098862
Rwpos5_15 in5 sp15 11140.846016
Rwpos5_16 in5 sp16 11140.846016
Rwpos5_17 in5 sp17 3183.098862
Rwpos5_18 in5 sp18 3183.098862
Rwpos5_19 in5 sp19 11140.846016
Rwpos5_20 in5 sp20 3183.098862
Rwpos5_21 in5 sp21 3183.098862
Rwpos5_22 in5 sp22 3183.098862
Rwpos5_23 in5 sp23 3183.098862
Rwpos5_24 in5 sp24 11140.846016
Rwpos5_25 in5 sp25 3183.098862
Rwpos5_26 in5 sp26 11140.846016
Rwpos5_27 in5 sp27 3183.098862
Rwpos5_28 in5 sp28 3183.098862
Rwpos5_29 in5 sp29 11140.846016
Rwpos5_30 in5 sp30 11140.846016
Rwpos5_31 in5 sp31 11140.846016
Rwpos5_32 in5 sp32 11140.846016
Rwpos5_33 in5 sp33 11140.846016
Rwpos5_34 in5 sp34 3183.098862
Rwpos5_35 in5 sp35 11140.846016
Rwpos5_36 in5 sp36 3183.098862
Rwpos5_37 in5 sp37 11140.846016
Rwpos5_38 in5 sp38 11140.846016
Rwpos5_39 in5 sp39 3183.098862
Rwpos5_40 in5 sp40 11140.846016
Rwpos5_41 in5 sp41 11140.846016
Rwpos5_42 in5 sp42 3183.098862
Rwpos5_43 in5 sp43 11140.846016
Rwpos5_44 in5 sp44 11140.846016
Rwpos5_45 in5 sp45 3183.098862
Rwpos5_46 in5 sp46 3183.098862
Rwpos5_47 in5 sp47 3183.098862
Rwpos5_48 in5 sp48 11140.846016
Rwpos5_49 in5 sp49 3183.098862
Rwpos5_50 in5 sp50 3183.098862
Rwpos5_51 in5 sp51 11140.846016
Rwpos5_52 in5 sp52 3183.098862
Rwpos5_53 in5 sp53 3183.098862
Rwpos5_54 in5 sp54 11140.846016
Rwpos5_55 in5 sp55 3183.098862
Rwpos5_56 in5 sp56 3183.098862
Rwpos5_57 in5 sp57 3183.098862
Rwpos5_58 in5 sp58 3183.098862
Rwpos5_59 in5 sp59 11140.846016
Rwpos5_60 in5 sp60 3183.098862
Rwpos5_61 in5 sp61 11140.846016
Rwpos5_62 in5 sp62 3183.098862
Rwpos5_63 in5 sp63 11140.846016
Rwpos5_64 in5 sp64 11140.846016
Rwpos5_65 in5 sp65 11140.846016
Rwpos5_66 in5 sp66 3183.098862
Rwpos5_67 in5 sp67 3183.098862
Rwpos5_68 in5 sp68 3183.098862
Rwpos5_69 in5 sp69 3183.098862
Rwpos5_70 in5 sp70 3183.098862
Rwpos5_71 in5 sp71 11140.846016
Rwpos5_72 in5 sp72 11140.846016
Rwpos5_73 in5 sp73 3183.098862
Rwpos5_74 in5 sp74 3183.098862
Rwpos5_75 in5 sp75 3183.098862
Rwpos5_76 in5 sp76 11140.846016
Rwpos5_77 in5 sp77 3183.098862
Rwpos5_78 in5 sp78 3183.098862
Rwpos5_79 in5 sp79 11140.846016
Rwpos5_80 in5 sp80 3183.098862
Rwpos5_81 in5 sp81 11140.846016
Rwpos5_82 in5 sp82 11140.846016
Rwpos5_83 in5 sp83 3183.098862
Rwpos5_84 in5 sp84 11140.846016
Rwpos5_85 in5 sp85 3183.098862
Rwpos5_86 in5 sp86 3183.098862
Rwpos5_87 in5 sp87 11140.846016
Rwpos5_88 in5 sp88 11140.846016
Rwpos5_89 in5 sp89 3183.098862
Rwpos5_90 in5 sp90 11140.846016
Rwpos5_91 in5 sp91 3183.098862
Rwpos5_92 in5 sp92 3183.098862
Rwpos5_93 in5 sp93 3183.098862
Rwpos5_94 in5 sp94 11140.846016
Rwpos5_95 in5 sp95 3183.098862
Rwpos5_96 in5 sp96 11140.846016
Rwpos5_97 in5 sp97 3183.098862
Rwpos5_98 in5 sp98 11140.846016
Rwpos5_99 in5 sp99 11140.846016
Rwpos5_100 in5 sp100 3183.098862
Rwpos6_1 in6 sp1 11140.846016
Rwpos6_2 in6 sp2 11140.846016
Rwpos6_3 in6 sp3 3183.098862
Rwpos6_4 in6 sp4 3183.098862
Rwpos6_5 in6 sp5 3183.098862
Rwpos6_6 in6 sp6 11140.846016
Rwpos6_7 in6 sp7 3183.098862
Rwpos6_8 in6 sp8 11140.846016
Rwpos6_9 in6 sp9 11140.846016
Rwpos6_10 in6 sp10 11140.846016
Rwpos6_11 in6 sp11 3183.098862
Rwpos6_12 in6 sp12 11140.846016
Rwpos6_13 in6 sp13 3183.098862
Rwpos6_14 in6 sp14 3183.098862
Rwpos6_15 in6 sp15 11140.846016
Rwpos6_16 in6 sp16 3183.098862
Rwpos6_17 in6 sp17 3183.098862
Rwpos6_18 in6 sp18 3183.098862
Rwpos6_19 in6 sp19 3183.098862
Rwpos6_20 in6 sp20 3183.098862
Rwpos6_21 in6 sp21 3183.098862
Rwpos6_22 in6 sp22 11140.846016
Rwpos6_23 in6 sp23 11140.846016
Rwpos6_24 in6 sp24 11140.846016
Rwpos6_25 in6 sp25 3183.098862
Rwpos6_26 in6 sp26 11140.846016
Rwpos6_27 in6 sp27 3183.098862
Rwpos6_28 in6 sp28 11140.846016
Rwpos6_29 in6 sp29 3183.098862
Rwpos6_30 in6 sp30 3183.098862
Rwpos6_31 in6 sp31 3183.098862
Rwpos6_32 in6 sp32 11140.846016
Rwpos6_33 in6 sp33 3183.098862
Rwpos6_34 in6 sp34 11140.846016
Rwpos6_35 in6 sp35 3183.098862
Rwpos6_36 in6 sp36 3183.098862
Rwpos6_37 in6 sp37 3183.098862
Rwpos6_38 in6 sp38 3183.098862
Rwpos6_39 in6 sp39 3183.098862
Rwpos6_40 in6 sp40 3183.098862
Rwpos6_41 in6 sp41 11140.846016
Rwpos6_42 in6 sp42 3183.098862
Rwpos6_43 in6 sp43 3183.098862
Rwpos6_44 in6 sp44 11140.846016
Rwpos6_45 in6 sp45 11140.846016
Rwpos6_46 in6 sp46 11140.846016
Rwpos6_47 in6 sp47 11140.846016
Rwpos6_48 in6 sp48 3183.098862
Rwpos6_49 in6 sp49 11140.846016
Rwpos6_50 in6 sp50 11140.846016
Rwpos6_51 in6 sp51 3183.098862
Rwpos6_52 in6 sp52 3183.098862
Rwpos6_53 in6 sp53 3183.098862
Rwpos6_54 in6 sp54 3183.098862
Rwpos6_55 in6 sp55 3183.098862
Rwpos6_56 in6 sp56 3183.098862
Rwpos6_57 in6 sp57 11140.846016
Rwpos6_58 in6 sp58 3183.098862
Rwpos6_59 in6 sp59 11140.846016
Rwpos6_60 in6 sp60 11140.846016
Rwpos6_61 in6 sp61 3183.098862
Rwpos6_62 in6 sp62 3183.098862
Rwpos6_63 in6 sp63 3183.098862
Rwpos6_64 in6 sp64 11140.846016
Rwpos6_65 in6 sp65 3183.098862
Rwpos6_66 in6 sp66 3183.098862
Rwpos6_67 in6 sp67 3183.098862
Rwpos6_68 in6 sp68 11140.846016
Rwpos6_69 in6 sp69 11140.846016
Rwpos6_70 in6 sp70 3183.098862
Rwpos6_71 in6 sp71 11140.846016
Rwpos6_72 in6 sp72 3183.098862
Rwpos6_73 in6 sp73 3183.098862
Rwpos6_74 in6 sp74 11140.846016
Rwpos6_75 in6 sp75 3183.098862
Rwpos6_76 in6 sp76 11140.846016
Rwpos6_77 in6 sp77 11140.846016
Rwpos6_78 in6 sp78 3183.098862
Rwpos6_79 in6 sp79 3183.098862
Rwpos6_80 in6 sp80 3183.098862
Rwpos6_81 in6 sp81 3183.098862
Rwpos6_82 in6 sp82 11140.846016
Rwpos6_83 in6 sp83 3183.098862
Rwpos6_84 in6 sp84 3183.098862
Rwpos6_85 in6 sp85 11140.846016
Rwpos6_86 in6 sp86 3183.098862
Rwpos6_87 in6 sp87 11140.846016
Rwpos6_88 in6 sp88 3183.098862
Rwpos6_89 in6 sp89 11140.846016
Rwpos6_90 in6 sp90 3183.098862
Rwpos6_91 in6 sp91 3183.098862
Rwpos6_92 in6 sp92 3183.098862
Rwpos6_93 in6 sp93 3183.098862
Rwpos6_94 in6 sp94 3183.098862
Rwpos6_95 in6 sp95 3183.098862
Rwpos6_96 in6 sp96 11140.846016
Rwpos6_97 in6 sp97 11140.846016
Rwpos6_98 in6 sp98 11140.846016
Rwpos6_99 in6 sp99 11140.846016
Rwpos6_100 in6 sp100 3183.098862
Rwpos7_1 in7 sp1 3183.098862
Rwpos7_2 in7 sp2 3183.098862
Rwpos7_3 in7 sp3 11140.846016
Rwpos7_4 in7 sp4 3183.098862
Rwpos7_5 in7 sp5 11140.846016
Rwpos7_6 in7 sp6 11140.846016
Rwpos7_7 in7 sp7 3183.098862
Rwpos7_8 in7 sp8 3183.098862
Rwpos7_9 in7 sp9 3183.098862
Rwpos7_10 in7 sp10 11140.846016
Rwpos7_11 in7 sp11 3183.098862
Rwpos7_12 in7 sp12 3183.098862
Rwpos7_13 in7 sp13 11140.846016
Rwpos7_14 in7 sp14 11140.846016
Rwpos7_15 in7 sp15 11140.846016
Rwpos7_16 in7 sp16 3183.098862
Rwpos7_17 in7 sp17 11140.846016
Rwpos7_18 in7 sp18 3183.098862
Rwpos7_19 in7 sp19 3183.098862
Rwpos7_20 in7 sp20 11140.846016
Rwpos7_21 in7 sp21 11140.846016
Rwpos7_22 in7 sp22 11140.846016
Rwpos7_23 in7 sp23 11140.846016
Rwpos7_24 in7 sp24 3183.098862
Rwpos7_25 in7 sp25 11140.846016
Rwpos7_26 in7 sp26 11140.846016
Rwpos7_27 in7 sp27 3183.098862
Rwpos7_28 in7 sp28 3183.098862
Rwpos7_29 in7 sp29 11140.846016
Rwpos7_30 in7 sp30 3183.098862
Rwpos7_31 in7 sp31 3183.098862
Rwpos7_32 in7 sp32 11140.846016
Rwpos7_33 in7 sp33 3183.098862
Rwpos7_34 in7 sp34 3183.098862
Rwpos7_35 in7 sp35 3183.098862
Rwpos7_36 in7 sp36 11140.846016
Rwpos7_37 in7 sp37 3183.098862
Rwpos7_38 in7 sp38 3183.098862
Rwpos7_39 in7 sp39 11140.846016
Rwpos7_40 in7 sp40 3183.098862
Rwpos7_41 in7 sp41 11140.846016
Rwpos7_42 in7 sp42 11140.846016
Rwpos7_43 in7 sp43 11140.846016
Rwpos7_44 in7 sp44 11140.846016
Rwpos7_45 in7 sp45 3183.098862
Rwpos7_46 in7 sp46 11140.846016
Rwpos7_47 in7 sp47 3183.098862
Rwpos7_48 in7 sp48 11140.846016
Rwpos7_49 in7 sp49 11140.846016
Rwpos7_50 in7 sp50 11140.846016
Rwpos7_51 in7 sp51 11140.846016
Rwpos7_52 in7 sp52 3183.098862
Rwpos7_53 in7 sp53 11140.846016
Rwpos7_54 in7 sp54 11140.846016
Rwpos7_55 in7 sp55 11140.846016
Rwpos7_56 in7 sp56 11140.846016
Rwpos7_57 in7 sp57 3183.098862
Rwpos7_58 in7 sp58 3183.098862
Rwpos7_59 in7 sp59 11140.846016
Rwpos7_60 in7 sp60 11140.846016
Rwpos7_61 in7 sp61 3183.098862
Rwpos7_62 in7 sp62 11140.846016
Rwpos7_63 in7 sp63 3183.098862
Rwpos7_64 in7 sp64 3183.098862
Rwpos7_65 in7 sp65 3183.098862
Rwpos7_66 in7 sp66 3183.098862
Rwpos7_67 in7 sp67 11140.846016
Rwpos7_68 in7 sp68 3183.098862
Rwpos7_69 in7 sp69 3183.098862
Rwpos7_70 in7 sp70 11140.846016
Rwpos7_71 in7 sp71 11140.846016
Rwpos7_72 in7 sp72 11140.846016
Rwpos7_73 in7 sp73 3183.098862
Rwpos7_74 in7 sp74 11140.846016
Rwpos7_75 in7 sp75 11140.846016
Rwpos7_76 in7 sp76 11140.846016
Rwpos7_77 in7 sp77 11140.846016
Rwpos7_78 in7 sp78 11140.846016
Rwpos7_79 in7 sp79 11140.846016
Rwpos7_80 in7 sp80 3183.098862
Rwpos7_81 in7 sp81 11140.846016
Rwpos7_82 in7 sp82 3183.098862
Rwpos7_83 in7 sp83 11140.846016
Rwpos7_84 in7 sp84 3183.098862
Rwpos7_85 in7 sp85 3183.098862
Rwpos7_86 in7 sp86 11140.846016
Rwpos7_87 in7 sp87 11140.846016
Rwpos7_88 in7 sp88 11140.846016
Rwpos7_89 in7 sp89 3183.098862
Rwpos7_90 in7 sp90 11140.846016
Rwpos7_91 in7 sp91 3183.098862
Rwpos7_92 in7 sp92 3183.098862
Rwpos7_93 in7 sp93 11140.846016
Rwpos7_94 in7 sp94 11140.846016
Rwpos7_95 in7 sp95 3183.098862
Rwpos7_96 in7 sp96 3183.098862
Rwpos7_97 in7 sp97 3183.098862
Rwpos7_98 in7 sp98 3183.098862
Rwpos7_99 in7 sp99 11140.846016
Rwpos7_100 in7 sp100 3183.098862
Rwpos8_1 in8 sp1 3183.098862
Rwpos8_2 in8 sp2 11140.846016
Rwpos8_3 in8 sp3 11140.846016
Rwpos8_4 in8 sp4 3183.098862
Rwpos8_5 in8 sp5 11140.846016
Rwpos8_6 in8 sp6 11140.846016
Rwpos8_7 in8 sp7 11140.846016
Rwpos8_8 in8 sp8 11140.846016
Rwpos8_9 in8 sp9 3183.098862
Rwpos8_10 in8 sp10 3183.098862
Rwpos8_11 in8 sp11 11140.846016
Rwpos8_12 in8 sp12 3183.098862
Rwpos8_13 in8 sp13 11140.846016
Rwpos8_14 in8 sp14 3183.098862
Rwpos8_15 in8 sp15 11140.846016
Rwpos8_16 in8 sp16 3183.098862
Rwpos8_17 in8 sp17 11140.846016
Rwpos8_18 in8 sp18 11140.846016
Rwpos8_19 in8 sp19 3183.098862
Rwpos8_20 in8 sp20 11140.846016
Rwpos8_21 in8 sp21 3183.098862
Rwpos8_22 in8 sp22 11140.846016
Rwpos8_23 in8 sp23 3183.098862
Rwpos8_24 in8 sp24 11140.846016
Rwpos8_25 in8 sp25 11140.846016
Rwpos8_26 in8 sp26 3183.098862
Rwpos8_27 in8 sp27 11140.846016
Rwpos8_28 in8 sp28 3183.098862
Rwpos8_29 in8 sp29 3183.098862
Rwpos8_30 in8 sp30 11140.846016
Rwpos8_31 in8 sp31 11140.846016
Rwpos8_32 in8 sp32 3183.098862
Rwpos8_33 in8 sp33 3183.098862
Rwpos8_34 in8 sp34 3183.098862
Rwpos8_35 in8 sp35 11140.846016
Rwpos8_36 in8 sp36 3183.098862
Rwpos8_37 in8 sp37 11140.846016
Rwpos8_38 in8 sp38 3183.098862
Rwpos8_39 in8 sp39 3183.098862
Rwpos8_40 in8 sp40 11140.846016
Rwpos8_41 in8 sp41 3183.098862
Rwpos8_42 in8 sp42 3183.098862
Rwpos8_43 in8 sp43 3183.098862
Rwpos8_44 in8 sp44 11140.846016
Rwpos8_45 in8 sp45 3183.098862
Rwpos8_46 in8 sp46 3183.098862
Rwpos8_47 in8 sp47 3183.098862
Rwpos8_48 in8 sp48 3183.098862
Rwpos8_49 in8 sp49 11140.846016
Rwpos8_50 in8 sp50 3183.098862
Rwpos8_51 in8 sp51 11140.846016
Rwpos8_52 in8 sp52 11140.846016
Rwpos8_53 in8 sp53 3183.098862
Rwpos8_54 in8 sp54 11140.846016
Rwpos8_55 in8 sp55 11140.846016
Rwpos8_56 in8 sp56 3183.098862
Rwpos8_57 in8 sp57 11140.846016
Rwpos8_58 in8 sp58 11140.846016
Rwpos8_59 in8 sp59 11140.846016
Rwpos8_60 in8 sp60 11140.846016
Rwpos8_61 in8 sp61 3183.098862
Rwpos8_62 in8 sp62 3183.098862
Rwpos8_63 in8 sp63 3183.098862
Rwpos8_64 in8 sp64 3183.098862
Rwpos8_65 in8 sp65 11140.846016
Rwpos8_66 in8 sp66 3183.098862
Rwpos8_67 in8 sp67 11140.846016
Rwpos8_68 in8 sp68 3183.098862
Rwpos8_69 in8 sp69 3183.098862
Rwpos8_70 in8 sp70 3183.098862
Rwpos8_71 in8 sp71 11140.846016
Rwpos8_72 in8 sp72 11140.846016
Rwpos8_73 in8 sp73 3183.098862
Rwpos8_74 in8 sp74 11140.846016
Rwpos8_75 in8 sp75 11140.846016
Rwpos8_76 in8 sp76 11140.846016
Rwpos8_77 in8 sp77 3183.098862
Rwpos8_78 in8 sp78 3183.098862
Rwpos8_79 in8 sp79 11140.846016
Rwpos8_80 in8 sp80 11140.846016
Rwpos8_81 in8 sp81 11140.846016
Rwpos8_82 in8 sp82 3183.098862
Rwpos8_83 in8 sp83 3183.098862
Rwpos8_84 in8 sp84 11140.846016
Rwpos8_85 in8 sp85 11140.846016
Rwpos8_86 in8 sp86 11140.846016
Rwpos8_87 in8 sp87 11140.846016
Rwpos8_88 in8 sp88 3183.098862
Rwpos8_89 in8 sp89 3183.098862
Rwpos8_90 in8 sp90 11140.846016
Rwpos8_91 in8 sp91 11140.846016
Rwpos8_92 in8 sp92 3183.098862
Rwpos8_93 in8 sp93 11140.846016
Rwpos8_94 in8 sp94 3183.098862
Rwpos8_95 in8 sp95 3183.098862
Rwpos8_96 in8 sp96 11140.846016
Rwpos8_97 in8 sp97 11140.846016
Rwpos8_98 in8 sp98 11140.846016
Rwpos8_99 in8 sp99 11140.846016
Rwpos8_100 in8 sp100 11140.846016
Rwpos9_1 in9 sp1 11140.846016
Rwpos9_2 in9 sp2 11140.846016
Rwpos9_3 in9 sp3 11140.846016
Rwpos9_4 in9 sp4 3183.098862
Rwpos9_5 in9 sp5 11140.846016
Rwpos9_6 in9 sp6 3183.098862
Rwpos9_7 in9 sp7 11140.846016
Rwpos9_8 in9 sp8 11140.846016
Rwpos9_9 in9 sp9 3183.098862
Rwpos9_10 in9 sp10 11140.846016
Rwpos9_11 in9 sp11 11140.846016
Rwpos9_12 in9 sp12 11140.846016
Rwpos9_13 in9 sp13 11140.846016
Rwpos9_14 in9 sp14 11140.846016
Rwpos9_15 in9 sp15 11140.846016
Rwpos9_16 in9 sp16 3183.098862
Rwpos9_17 in9 sp17 3183.098862
Rwpos9_18 in9 sp18 3183.098862
Rwpos9_19 in9 sp19 11140.846016
Rwpos9_20 in9 sp20 11140.846016
Rwpos9_21 in9 sp21 3183.098862
Rwpos9_22 in9 sp22 11140.846016
Rwpos9_23 in9 sp23 11140.846016
Rwpos9_24 in9 sp24 3183.098862
Rwpos9_25 in9 sp25 3183.098862
Rwpos9_26 in9 sp26 3183.098862
Rwpos9_27 in9 sp27 3183.098862
Rwpos9_28 in9 sp28 11140.846016
Rwpos9_29 in9 sp29 3183.098862
Rwpos9_30 in9 sp30 11140.846016
Rwpos9_31 in9 sp31 3183.098862
Rwpos9_32 in9 sp32 11140.846016
Rwpos9_33 in9 sp33 3183.098862
Rwpos9_34 in9 sp34 11140.846016
Rwpos9_35 in9 sp35 11140.846016
Rwpos9_36 in9 sp36 11140.846016
Rwpos9_37 in9 sp37 3183.098862
Rwpos9_38 in9 sp38 11140.846016
Rwpos9_39 in9 sp39 3183.098862
Rwpos9_40 in9 sp40 3183.098862
Rwpos9_41 in9 sp41 3183.098862
Rwpos9_42 in9 sp42 11140.846016
Rwpos9_43 in9 sp43 11140.846016
Rwpos9_44 in9 sp44 3183.098862
Rwpos9_45 in9 sp45 11140.846016
Rwpos9_46 in9 sp46 11140.846016
Rwpos9_47 in9 sp47 3183.098862
Rwpos9_48 in9 sp48 11140.846016
Rwpos9_49 in9 sp49 11140.846016
Rwpos9_50 in9 sp50 11140.846016
Rwpos9_51 in9 sp51 11140.846016
Rwpos9_52 in9 sp52 3183.098862
Rwpos9_53 in9 sp53 3183.098862
Rwpos9_54 in9 sp54 11140.846016
Rwpos9_55 in9 sp55 11140.846016
Rwpos9_56 in9 sp56 3183.098862
Rwpos9_57 in9 sp57 11140.846016
Rwpos9_58 in9 sp58 3183.098862
Rwpos9_59 in9 sp59 11140.846016
Rwpos9_60 in9 sp60 11140.846016
Rwpos9_61 in9 sp61 3183.098862
Rwpos9_62 in9 sp62 11140.846016
Rwpos9_63 in9 sp63 3183.098862
Rwpos9_64 in9 sp64 3183.098862
Rwpos9_65 in9 sp65 3183.098862
Rwpos9_66 in9 sp66 11140.846016
Rwpos9_67 in9 sp67 3183.098862
Rwpos9_68 in9 sp68 11140.846016
Rwpos9_69 in9 sp69 3183.098862
Rwpos9_70 in9 sp70 11140.846016
Rwpos9_71 in9 sp71 11140.846016
Rwpos9_72 in9 sp72 11140.846016
Rwpos9_73 in9 sp73 11140.846016
Rwpos9_74 in9 sp74 3183.098862
Rwpos9_75 in9 sp75 3183.098862
Rwpos9_76 in9 sp76 11140.846016
Rwpos9_77 in9 sp77 3183.098862
Rwpos9_78 in9 sp78 11140.846016
Rwpos9_79 in9 sp79 3183.098862
Rwpos9_80 in9 sp80 11140.846016
Rwpos9_81 in9 sp81 11140.846016
Rwpos9_82 in9 sp82 3183.098862
Rwpos9_83 in9 sp83 3183.098862
Rwpos9_84 in9 sp84 11140.846016
Rwpos9_85 in9 sp85 3183.098862
Rwpos9_86 in9 sp86 11140.846016
Rwpos9_87 in9 sp87 11140.846016
Rwpos9_88 in9 sp88 3183.098862
Rwpos9_89 in9 sp89 3183.098862
Rwpos9_90 in9 sp90 11140.846016
Rwpos9_91 in9 sp91 3183.098862
Rwpos9_92 in9 sp92 3183.098862
Rwpos9_93 in9 sp93 11140.846016
Rwpos9_94 in9 sp94 3183.098862
Rwpos9_95 in9 sp95 3183.098862
Rwpos9_96 in9 sp96 11140.846016
Rwpos9_97 in9 sp97 11140.846016
Rwpos9_98 in9 sp98 3183.098862
Rwpos9_99 in9 sp99 11140.846016
Rwpos9_100 in9 sp100 3183.098862
Rwpos10_1 in10 sp1 11140.846016
Rwpos10_2 in10 sp2 11140.846016
Rwpos10_3 in10 sp3 11140.846016
Rwpos10_4 in10 sp4 3183.098862
Rwpos10_5 in10 sp5 11140.846016
Rwpos10_6 in10 sp6 11140.846016
Rwpos10_7 in10 sp7 11140.846016
Rwpos10_8 in10 sp8 11140.846016
Rwpos10_9 in10 sp9 3183.098862
Rwpos10_10 in10 sp10 3183.098862
Rwpos10_11 in10 sp11 3183.098862
Rwpos10_12 in10 sp12 11140.846016
Rwpos10_13 in10 sp13 3183.098862
Rwpos10_14 in10 sp14 11140.846016
Rwpos10_15 in10 sp15 11140.846016
Rwpos10_16 in10 sp16 11140.846016
Rwpos10_17 in10 sp17 11140.846016
Rwpos10_18 in10 sp18 11140.846016
Rwpos10_19 in10 sp19 11140.846016
Rwpos10_20 in10 sp20 11140.846016
Rwpos10_21 in10 sp21 3183.098862
Rwpos10_22 in10 sp22 3183.098862
Rwpos10_23 in10 sp23 3183.098862
Rwpos10_24 in10 sp24 3183.098862
Rwpos10_25 in10 sp25 11140.846016
Rwpos10_26 in10 sp26 3183.098862
Rwpos10_27 in10 sp27 11140.846016
Rwpos10_28 in10 sp28 11140.846016
Rwpos10_29 in10 sp29 3183.098862
Rwpos10_30 in10 sp30 11140.846016
Rwpos10_31 in10 sp31 11140.846016
Rwpos10_32 in10 sp32 11140.846016
Rwpos10_33 in10 sp33 11140.846016
Rwpos10_34 in10 sp34 3183.098862
Rwpos10_35 in10 sp35 11140.846016
Rwpos10_36 in10 sp36 3183.098862
Rwpos10_37 in10 sp37 3183.098862
Rwpos10_38 in10 sp38 3183.098862
Rwpos10_39 in10 sp39 3183.098862
Rwpos10_40 in10 sp40 11140.846016
Rwpos10_41 in10 sp41 11140.846016
Rwpos10_42 in10 sp42 11140.846016
Rwpos10_43 in10 sp43 3183.098862
Rwpos10_44 in10 sp44 3183.098862
Rwpos10_45 in10 sp45 11140.846016
Rwpos10_46 in10 sp46 3183.098862
Rwpos10_47 in10 sp47 3183.098862
Rwpos10_48 in10 sp48 3183.098862
Rwpos10_49 in10 sp49 11140.846016
Rwpos10_50 in10 sp50 3183.098862
Rwpos10_51 in10 sp51 11140.846016
Rwpos10_52 in10 sp52 3183.098862
Rwpos10_53 in10 sp53 11140.846016
Rwpos10_54 in10 sp54 11140.846016
Rwpos10_55 in10 sp55 11140.846016
Rwpos10_56 in10 sp56 11140.846016
Rwpos10_57 in10 sp57 11140.846016
Rwpos10_58 in10 sp58 11140.846016
Rwpos10_59 in10 sp59 3183.098862
Rwpos10_60 in10 sp60 3183.098862
Rwpos10_61 in10 sp61 11140.846016
Rwpos10_62 in10 sp62 3183.098862
Rwpos10_63 in10 sp63 3183.098862
Rwpos10_64 in10 sp64 11140.846016
Rwpos10_65 in10 sp65 11140.846016
Rwpos10_66 in10 sp66 11140.846016
Rwpos10_67 in10 sp67 11140.846016
Rwpos10_68 in10 sp68 11140.846016
Rwpos10_69 in10 sp69 3183.098862
Rwpos10_70 in10 sp70 11140.846016
Rwpos10_71 in10 sp71 11140.846016
Rwpos10_72 in10 sp72 11140.846016
Rwpos10_73 in10 sp73 11140.846016
Rwpos10_74 in10 sp74 3183.098862
Rwpos10_75 in10 sp75 3183.098862
Rwpos10_76 in10 sp76 3183.098862
Rwpos10_77 in10 sp77 11140.846016
Rwpos10_78 in10 sp78 11140.846016
Rwpos10_79 in10 sp79 3183.098862
Rwpos10_80 in10 sp80 11140.846016
Rwpos10_81 in10 sp81 11140.846016
Rwpos10_82 in10 sp82 11140.846016
Rwpos10_83 in10 sp83 3183.098862
Rwpos10_84 in10 sp84 11140.846016
Rwpos10_85 in10 sp85 3183.098862
Rwpos10_86 in10 sp86 3183.098862
Rwpos10_87 in10 sp87 11140.846016
Rwpos10_88 in10 sp88 3183.098862
Rwpos10_89 in10 sp89 11140.846016
Rwpos10_90 in10 sp90 11140.846016
Rwpos10_91 in10 sp91 3183.098862
Rwpos10_92 in10 sp92 3183.098862
Rwpos10_93 in10 sp93 11140.846016
Rwpos10_94 in10 sp94 11140.846016
Rwpos10_95 in10 sp95 11140.846016
Rwpos10_96 in10 sp96 3183.098862
Rwpos10_97 in10 sp97 3183.098862
Rwpos10_98 in10 sp98 3183.098862
Rwpos10_99 in10 sp99 11140.846016
Rwpos10_100 in10 sp100 3183.098862
Rwpos11_1 in11 sp1 3183.098862
Rwpos11_2 in11 sp2 3183.098862
Rwpos11_3 in11 sp3 3183.098862
Rwpos11_4 in11 sp4 3183.098862
Rwpos11_5 in11 sp5 11140.846016
Rwpos11_6 in11 sp6 11140.846016
Rwpos11_7 in11 sp7 11140.846016
Rwpos11_8 in11 sp8 11140.846016
Rwpos11_9 in11 sp9 3183.098862
Rwpos11_10 in11 sp10 3183.098862
Rwpos11_11 in11 sp11 3183.098862
Rwpos11_12 in11 sp12 3183.098862
Rwpos11_13 in11 sp13 3183.098862
Rwpos11_14 in11 sp14 3183.098862
Rwpos11_15 in11 sp15 11140.846016
Rwpos11_16 in11 sp16 11140.846016
Rwpos11_17 in11 sp17 11140.846016
Rwpos11_18 in11 sp18 3183.098862
Rwpos11_19 in11 sp19 3183.098862
Rwpos11_20 in11 sp20 3183.098862
Rwpos11_21 in11 sp21 11140.846016
Rwpos11_22 in11 sp22 3183.098862
Rwpos11_23 in11 sp23 11140.846016
Rwpos11_24 in11 sp24 11140.846016
Rwpos11_25 in11 sp25 3183.098862
Rwpos11_26 in11 sp26 3183.098862
Rwpos11_27 in11 sp27 3183.098862
Rwpos11_28 in11 sp28 3183.098862
Rwpos11_29 in11 sp29 3183.098862
Rwpos11_30 in11 sp30 3183.098862
Rwpos11_31 in11 sp31 3183.098862
Rwpos11_32 in11 sp32 3183.098862
Rwpos11_33 in11 sp33 11140.846016
Rwpos11_34 in11 sp34 11140.846016
Rwpos11_35 in11 sp35 11140.846016
Rwpos11_36 in11 sp36 3183.098862
Rwpos11_37 in11 sp37 3183.098862
Rwpos11_38 in11 sp38 11140.846016
Rwpos11_39 in11 sp39 3183.098862
Rwpos11_40 in11 sp40 11140.846016
Rwpos11_41 in11 sp41 11140.846016
Rwpos11_42 in11 sp42 3183.098862
Rwpos11_43 in11 sp43 3183.098862
Rwpos11_44 in11 sp44 11140.846016
Rwpos11_45 in11 sp45 11140.846016
Rwpos11_46 in11 sp46 3183.098862
Rwpos11_47 in11 sp47 3183.098862
Rwpos11_48 in11 sp48 11140.846016
Rwpos11_49 in11 sp49 11140.846016
Rwpos11_50 in11 sp50 11140.846016
Rwpos11_51 in11 sp51 11140.846016
Rwpos11_52 in11 sp52 3183.098862
Rwpos11_53 in11 sp53 11140.846016
Rwpos11_54 in11 sp54 11140.846016
Rwpos11_55 in11 sp55 11140.846016
Rwpos11_56 in11 sp56 3183.098862
Rwpos11_57 in11 sp57 3183.098862
Rwpos11_58 in11 sp58 11140.846016
Rwpos11_59 in11 sp59 3183.098862
Rwpos11_60 in11 sp60 11140.846016
Rwpos11_61 in11 sp61 3183.098862
Rwpos11_62 in11 sp62 11140.846016
Rwpos11_63 in11 sp63 3183.098862
Rwpos11_64 in11 sp64 11140.846016
Rwpos11_65 in11 sp65 11140.846016
Rwpos11_66 in11 sp66 3183.098862
Rwpos11_67 in11 sp67 3183.098862
Rwpos11_68 in11 sp68 3183.098862
Rwpos11_69 in11 sp69 3183.098862
Rwpos11_70 in11 sp70 3183.098862
Rwpos11_71 in11 sp71 11140.846016
Rwpos11_72 in11 sp72 11140.846016
Rwpos11_73 in11 sp73 3183.098862
Rwpos11_74 in11 sp74 3183.098862
Rwpos11_75 in11 sp75 3183.098862
Rwpos11_76 in11 sp76 3183.098862
Rwpos11_77 in11 sp77 3183.098862
Rwpos11_78 in11 sp78 3183.098862
Rwpos11_79 in11 sp79 11140.846016
Rwpos11_80 in11 sp80 11140.846016
Rwpos11_81 in11 sp81 3183.098862
Rwpos11_82 in11 sp82 11140.846016
Rwpos11_83 in11 sp83 11140.846016
Rwpos11_84 in11 sp84 11140.846016
Rwpos11_85 in11 sp85 3183.098862
Rwpos11_86 in11 sp86 11140.846016
Rwpos11_87 in11 sp87 3183.098862
Rwpos11_88 in11 sp88 3183.098862
Rwpos11_89 in11 sp89 3183.098862
Rwpos11_90 in11 sp90 3183.098862
Rwpos11_91 in11 sp91 3183.098862
Rwpos11_92 in11 sp92 3183.098862
Rwpos11_93 in11 sp93 3183.098862
Rwpos11_94 in11 sp94 11140.846016
Rwpos11_95 in11 sp95 11140.846016
Rwpos11_96 in11 sp96 3183.098862
Rwpos11_97 in11 sp97 3183.098862
Rwpos11_98 in11 sp98 11140.846016
Rwpos11_99 in11 sp99 3183.098862
Rwpos11_100 in11 sp100 3183.098862
Rwpos12_1 in12 sp1 11140.846016
Rwpos12_2 in12 sp2 3183.098862
Rwpos12_3 in12 sp3 3183.098862
Rwpos12_4 in12 sp4 11140.846016
Rwpos12_5 in12 sp5 3183.098862
Rwpos12_6 in12 sp6 3183.098862
Rwpos12_7 in12 sp7 3183.098862
Rwpos12_8 in12 sp8 11140.846016
Rwpos12_9 in12 sp9 3183.098862
Rwpos12_10 in12 sp10 11140.846016
Rwpos12_11 in12 sp11 3183.098862
Rwpos12_12 in12 sp12 3183.098862
Rwpos12_13 in12 sp13 11140.846016
Rwpos12_14 in12 sp14 11140.846016
Rwpos12_15 in12 sp15 3183.098862
Rwpos12_16 in12 sp16 3183.098862
Rwpos12_17 in12 sp17 3183.098862
Rwpos12_18 in12 sp18 3183.098862
Rwpos12_19 in12 sp19 3183.098862
Rwpos12_20 in12 sp20 11140.846016
Rwpos12_21 in12 sp21 11140.846016
Rwpos12_22 in12 sp22 3183.098862
Rwpos12_23 in12 sp23 3183.098862
Rwpos12_24 in12 sp24 3183.098862
Rwpos12_25 in12 sp25 11140.846016
Rwpos12_26 in12 sp26 11140.846016
Rwpos12_27 in12 sp27 3183.098862
Rwpos12_28 in12 sp28 3183.098862
Rwpos12_29 in12 sp29 11140.846016
Rwpos12_30 in12 sp30 11140.846016
Rwpos12_31 in12 sp31 11140.846016
Rwpos12_32 in12 sp32 3183.098862
Rwpos12_33 in12 sp33 3183.098862
Rwpos12_34 in12 sp34 3183.098862
Rwpos12_35 in12 sp35 3183.098862
Rwpos12_36 in12 sp36 11140.846016
Rwpos12_37 in12 sp37 3183.098862
Rwpos12_38 in12 sp38 11140.846016
Rwpos12_39 in12 sp39 3183.098862
Rwpos12_40 in12 sp40 3183.098862
Rwpos12_41 in12 sp41 3183.098862
Rwpos12_42 in12 sp42 11140.846016
Rwpos12_43 in12 sp43 3183.098862
Rwpos12_44 in12 sp44 3183.098862
Rwpos12_45 in12 sp45 3183.098862
Rwpos12_46 in12 sp46 3183.098862
Rwpos12_47 in12 sp47 11140.846016
Rwpos12_48 in12 sp48 3183.098862
Rwpos12_49 in12 sp49 3183.098862
Rwpos12_50 in12 sp50 3183.098862
Rwpos12_51 in12 sp51 11140.846016
Rwpos12_52 in12 sp52 11140.846016
Rwpos12_53 in12 sp53 3183.098862
Rwpos12_54 in12 sp54 3183.098862
Rwpos12_55 in12 sp55 3183.098862
Rwpos12_56 in12 sp56 11140.846016
Rwpos12_57 in12 sp57 11140.846016
Rwpos12_58 in12 sp58 11140.846016
Rwpos12_59 in12 sp59 3183.098862
Rwpos12_60 in12 sp60 3183.098862
Rwpos12_61 in12 sp61 3183.098862
Rwpos12_62 in12 sp62 11140.846016
Rwpos12_63 in12 sp63 11140.846016
Rwpos12_64 in12 sp64 11140.846016
Rwpos12_65 in12 sp65 11140.846016
Rwpos12_66 in12 sp66 11140.846016
Rwpos12_67 in12 sp67 3183.098862
Rwpos12_68 in12 sp68 3183.098862
Rwpos12_69 in12 sp69 11140.846016
Rwpos12_70 in12 sp70 3183.098862
Rwpos12_71 in12 sp71 11140.846016
Rwpos12_72 in12 sp72 3183.098862
Rwpos12_73 in12 sp73 3183.098862
Rwpos12_74 in12 sp74 11140.846016
Rwpos12_75 in12 sp75 3183.098862
Rwpos12_76 in12 sp76 3183.098862
Rwpos12_77 in12 sp77 3183.098862
Rwpos12_78 in12 sp78 3183.098862
Rwpos12_79 in12 sp79 3183.098862
Rwpos12_80 in12 sp80 3183.098862
Rwpos12_81 in12 sp81 11140.846016
Rwpos12_82 in12 sp82 3183.098862
Rwpos12_83 in12 sp83 11140.846016
Rwpos12_84 in12 sp84 11140.846016
Rwpos12_85 in12 sp85 3183.098862
Rwpos12_86 in12 sp86 3183.098862
Rwpos12_87 in12 sp87 11140.846016
Rwpos12_88 in12 sp88 11140.846016
Rwpos12_89 in12 sp89 11140.846016
Rwpos12_90 in12 sp90 11140.846016
Rwpos12_91 in12 sp91 3183.098862
Rwpos12_92 in12 sp92 3183.098862
Rwpos12_93 in12 sp93 3183.098862
Rwpos12_94 in12 sp94 11140.846016
Rwpos12_95 in12 sp95 3183.098862
Rwpos12_96 in12 sp96 3183.098862
Rwpos12_97 in12 sp97 11140.846016
Rwpos12_98 in12 sp98 3183.098862
Rwpos12_99 in12 sp99 11140.846016
Rwpos12_100 in12 sp100 11140.846016
Rwpos13_1 in13 sp1 3183.098862
Rwpos13_2 in13 sp2 3183.098862
Rwpos13_3 in13 sp3 3183.098862
Rwpos13_4 in13 sp4 3183.098862
Rwpos13_5 in13 sp5 11140.846016
Rwpos13_6 in13 sp6 3183.098862
Rwpos13_7 in13 sp7 3183.098862
Rwpos13_8 in13 sp8 3183.098862
Rwpos13_9 in13 sp9 3183.098862
Rwpos13_10 in13 sp10 11140.846016
Rwpos13_11 in13 sp11 11140.846016
Rwpos13_12 in13 sp12 3183.098862
Rwpos13_13 in13 sp13 3183.098862
Rwpos13_14 in13 sp14 3183.098862
Rwpos13_15 in13 sp15 11140.846016
Rwpos13_16 in13 sp16 3183.098862
Rwpos13_17 in13 sp17 11140.846016
Rwpos13_18 in13 sp18 11140.846016
Rwpos13_19 in13 sp19 11140.846016
Rwpos13_20 in13 sp20 11140.846016
Rwpos13_21 in13 sp21 3183.098862
Rwpos13_22 in13 sp22 11140.846016
Rwpos13_23 in13 sp23 3183.098862
Rwpos13_24 in13 sp24 11140.846016
Rwpos13_25 in13 sp25 11140.846016
Rwpos13_26 in13 sp26 11140.846016
Rwpos13_27 in13 sp27 3183.098862
Rwpos13_28 in13 sp28 3183.098862
Rwpos13_29 in13 sp29 11140.846016
Rwpos13_30 in13 sp30 3183.098862
Rwpos13_31 in13 sp31 11140.846016
Rwpos13_32 in13 sp32 11140.846016
Rwpos13_33 in13 sp33 3183.098862
Rwpos13_34 in13 sp34 3183.098862
Rwpos13_35 in13 sp35 3183.098862
Rwpos13_36 in13 sp36 11140.846016
Rwpos13_37 in13 sp37 11140.846016
Rwpos13_38 in13 sp38 11140.846016
Rwpos13_39 in13 sp39 11140.846016
Rwpos13_40 in13 sp40 3183.098862
Rwpos13_41 in13 sp41 11140.846016
Rwpos13_42 in13 sp42 3183.098862
Rwpos13_43 in13 sp43 11140.846016
Rwpos13_44 in13 sp44 11140.846016
Rwpos13_45 in13 sp45 3183.098862
Rwpos13_46 in13 sp46 3183.098862
Rwpos13_47 in13 sp47 3183.098862
Rwpos13_48 in13 sp48 3183.098862
Rwpos13_49 in13 sp49 11140.846016
Rwpos13_50 in13 sp50 11140.846016
Rwpos13_51 in13 sp51 11140.846016
Rwpos13_52 in13 sp52 11140.846016
Rwpos13_53 in13 sp53 3183.098862
Rwpos13_54 in13 sp54 11140.846016
Rwpos13_55 in13 sp55 11140.846016
Rwpos13_56 in13 sp56 11140.846016
Rwpos13_57 in13 sp57 3183.098862
Rwpos13_58 in13 sp58 3183.098862
Rwpos13_59 in13 sp59 11140.846016
Rwpos13_60 in13 sp60 3183.098862
Rwpos13_61 in13 sp61 11140.846016
Rwpos13_62 in13 sp62 3183.098862
Rwpos13_63 in13 sp63 3183.098862
Rwpos13_64 in13 sp64 3183.098862
Rwpos13_65 in13 sp65 11140.846016
Rwpos13_66 in13 sp66 11140.846016
Rwpos13_67 in13 sp67 11140.846016
Rwpos13_68 in13 sp68 3183.098862
Rwpos13_69 in13 sp69 11140.846016
Rwpos13_70 in13 sp70 11140.846016
Rwpos13_71 in13 sp71 3183.098862
Rwpos13_72 in13 sp72 11140.846016
Rwpos13_73 in13 sp73 11140.846016
Rwpos13_74 in13 sp74 3183.098862
Rwpos13_75 in13 sp75 3183.098862
Rwpos13_76 in13 sp76 11140.846016
Rwpos13_77 in13 sp77 11140.846016
Rwpos13_78 in13 sp78 3183.098862
Rwpos13_79 in13 sp79 11140.846016
Rwpos13_80 in13 sp80 11140.846016
Rwpos13_81 in13 sp81 3183.098862
Rwpos13_82 in13 sp82 3183.098862
Rwpos13_83 in13 sp83 11140.846016
Rwpos13_84 in13 sp84 11140.846016
Rwpos13_85 in13 sp85 11140.846016
Rwpos13_86 in13 sp86 11140.846016
Rwpos13_87 in13 sp87 11140.846016
Rwpos13_88 in13 sp88 3183.098862
Rwpos13_89 in13 sp89 3183.098862
Rwpos13_90 in13 sp90 3183.098862
Rwpos13_91 in13 sp91 11140.846016
Rwpos13_92 in13 sp92 11140.846016
Rwpos13_93 in13 sp93 3183.098862
Rwpos13_94 in13 sp94 3183.098862
Rwpos13_95 in13 sp95 11140.846016
Rwpos13_96 in13 sp96 3183.098862
Rwpos13_97 in13 sp97 3183.098862
Rwpos13_98 in13 sp98 3183.098862
Rwpos13_99 in13 sp99 11140.846016
Rwpos13_100 in13 sp100 3183.098862
Rwpos14_1 in14 sp1 11140.846016
Rwpos14_2 in14 sp2 11140.846016
Rwpos14_3 in14 sp3 11140.846016
Rwpos14_4 in14 sp4 3183.098862
Rwpos14_5 in14 sp5 11140.846016
Rwpos14_6 in14 sp6 11140.846016
Rwpos14_7 in14 sp7 3183.098862
Rwpos14_8 in14 sp8 3183.098862
Rwpos14_9 in14 sp9 11140.846016
Rwpos14_10 in14 sp10 3183.098862
Rwpos14_11 in14 sp11 3183.098862
Rwpos14_12 in14 sp12 3183.098862
Rwpos14_13 in14 sp13 3183.098862
Rwpos14_14 in14 sp14 3183.098862
Rwpos14_15 in14 sp15 11140.846016
Rwpos14_16 in14 sp16 11140.846016
Rwpos14_17 in14 sp17 3183.098862
Rwpos14_18 in14 sp18 3183.098862
Rwpos14_19 in14 sp19 3183.098862
Rwpos14_20 in14 sp20 11140.846016
Rwpos14_21 in14 sp21 3183.098862
Rwpos14_22 in14 sp22 3183.098862
Rwpos14_23 in14 sp23 3183.098862
Rwpos14_24 in14 sp24 3183.098862
Rwpos14_25 in14 sp25 3183.098862
Rwpos14_26 in14 sp26 3183.098862
Rwpos14_27 in14 sp27 11140.846016
Rwpos14_28 in14 sp28 11140.846016
Rwpos14_29 in14 sp29 11140.846016
Rwpos14_30 in14 sp30 3183.098862
Rwpos14_31 in14 sp31 3183.098862
Rwpos14_32 in14 sp32 3183.098862
Rwpos14_33 in14 sp33 3183.098862
Rwpos14_34 in14 sp34 11140.846016
Rwpos14_35 in14 sp35 11140.846016
Rwpos14_36 in14 sp36 11140.846016
Rwpos14_37 in14 sp37 11140.846016
Rwpos14_38 in14 sp38 3183.098862
Rwpos14_39 in14 sp39 11140.846016
Rwpos14_40 in14 sp40 3183.098862
Rwpos14_41 in14 sp41 3183.098862
Rwpos14_42 in14 sp42 11140.846016
Rwpos14_43 in14 sp43 11140.846016
Rwpos14_44 in14 sp44 3183.098862
Rwpos14_45 in14 sp45 11140.846016
Rwpos14_46 in14 sp46 11140.846016
Rwpos14_47 in14 sp47 11140.846016
Rwpos14_48 in14 sp48 3183.098862
Rwpos14_49 in14 sp49 11140.846016
Rwpos14_50 in14 sp50 3183.098862
Rwpos14_51 in14 sp51 11140.846016
Rwpos14_52 in14 sp52 3183.098862
Rwpos14_53 in14 sp53 3183.098862
Rwpos14_54 in14 sp54 11140.846016
Rwpos14_55 in14 sp55 11140.846016
Rwpos14_56 in14 sp56 11140.846016
Rwpos14_57 in14 sp57 11140.846016
Rwpos14_58 in14 sp58 3183.098862
Rwpos14_59 in14 sp59 3183.098862
Rwpos14_60 in14 sp60 11140.846016
Rwpos14_61 in14 sp61 11140.846016
Rwpos14_62 in14 sp62 3183.098862
Rwpos14_63 in14 sp63 3183.098862
Rwpos14_64 in14 sp64 3183.098862
Rwpos14_65 in14 sp65 3183.098862
Rwpos14_66 in14 sp66 3183.098862
Rwpos14_67 in14 sp67 11140.846016
Rwpos14_68 in14 sp68 11140.846016
Rwpos14_69 in14 sp69 3183.098862
Rwpos14_70 in14 sp70 11140.846016
Rwpos14_71 in14 sp71 11140.846016
Rwpos14_72 in14 sp72 3183.098862
Rwpos14_73 in14 sp73 3183.098862
Rwpos14_74 in14 sp74 3183.098862
Rwpos14_75 in14 sp75 3183.098862
Rwpos14_76 in14 sp76 11140.846016
Rwpos14_77 in14 sp77 3183.098862
Rwpos14_78 in14 sp78 11140.846016
Rwpos14_79 in14 sp79 3183.098862
Rwpos14_80 in14 sp80 11140.846016
Rwpos14_81 in14 sp81 11140.846016
Rwpos14_82 in14 sp82 11140.846016
Rwpos14_83 in14 sp83 11140.846016
Rwpos14_84 in14 sp84 3183.098862
Rwpos14_85 in14 sp85 3183.098862
Rwpos14_86 in14 sp86 11140.846016
Rwpos14_87 in14 sp87 11140.846016
Rwpos14_88 in14 sp88 11140.846016
Rwpos14_89 in14 sp89 11140.846016
Rwpos14_90 in14 sp90 3183.098862
Rwpos14_91 in14 sp91 3183.098862
Rwpos14_92 in14 sp92 11140.846016
Rwpos14_93 in14 sp93 11140.846016
Rwpos14_94 in14 sp94 3183.098862
Rwpos14_95 in14 sp95 3183.098862
Rwpos14_96 in14 sp96 3183.098862
Rwpos14_97 in14 sp97 11140.846016
Rwpos14_98 in14 sp98 11140.846016
Rwpos14_99 in14 sp99 11140.846016
Rwpos14_100 in14 sp100 11140.846016
Rwpos15_1 in15 sp1 11140.846016
Rwpos15_2 in15 sp2 11140.846016
Rwpos15_3 in15 sp3 3183.098862
Rwpos15_4 in15 sp4 3183.098862
Rwpos15_5 in15 sp5 3183.098862
Rwpos15_6 in15 sp6 11140.846016
Rwpos15_7 in15 sp7 11140.846016
Rwpos15_8 in15 sp8 11140.846016
Rwpos15_9 in15 sp9 11140.846016
Rwpos15_10 in15 sp10 3183.098862
Rwpos15_11 in15 sp11 11140.846016
Rwpos15_12 in15 sp12 11140.846016
Rwpos15_13 in15 sp13 11140.846016
Rwpos15_14 in15 sp14 3183.098862
Rwpos15_15 in15 sp15 3183.098862
Rwpos15_16 in15 sp16 11140.846016
Rwpos15_17 in15 sp17 11140.846016
Rwpos15_18 in15 sp18 11140.846016
Rwpos15_19 in15 sp19 11140.846016
Rwpos15_20 in15 sp20 11140.846016
Rwpos15_21 in15 sp21 3183.098862
Rwpos15_22 in15 sp22 3183.098862
Rwpos15_23 in15 sp23 11140.846016
Rwpos15_24 in15 sp24 3183.098862
Rwpos15_25 in15 sp25 11140.846016
Rwpos15_26 in15 sp26 11140.846016
Rwpos15_27 in15 sp27 11140.846016
Rwpos15_28 in15 sp28 3183.098862
Rwpos15_29 in15 sp29 11140.846016
Rwpos15_30 in15 sp30 3183.098862
Rwpos15_31 in15 sp31 3183.098862
Rwpos15_32 in15 sp32 3183.098862
Rwpos15_33 in15 sp33 3183.098862
Rwpos15_34 in15 sp34 3183.098862
Rwpos15_35 in15 sp35 3183.098862
Rwpos15_36 in15 sp36 11140.846016
Rwpos15_37 in15 sp37 3183.098862
Rwpos15_38 in15 sp38 3183.098862
Rwpos15_39 in15 sp39 3183.098862
Rwpos15_40 in15 sp40 11140.846016
Rwpos15_41 in15 sp41 11140.846016
Rwpos15_42 in15 sp42 3183.098862
Rwpos15_43 in15 sp43 11140.846016
Rwpos15_44 in15 sp44 11140.846016
Rwpos15_45 in15 sp45 11140.846016
Rwpos15_46 in15 sp46 11140.846016
Rwpos15_47 in15 sp47 11140.846016
Rwpos15_48 in15 sp48 11140.846016
Rwpos15_49 in15 sp49 3183.098862
Rwpos15_50 in15 sp50 11140.846016
Rwpos15_51 in15 sp51 3183.098862
Rwpos15_52 in15 sp52 3183.098862
Rwpos15_53 in15 sp53 11140.846016
Rwpos15_54 in15 sp54 11140.846016
Rwpos15_55 in15 sp55 11140.846016
Rwpos15_56 in15 sp56 3183.098862
Rwpos15_57 in15 sp57 3183.098862
Rwpos15_58 in15 sp58 3183.098862
Rwpos15_59 in15 sp59 3183.098862
Rwpos15_60 in15 sp60 11140.846016
Rwpos15_61 in15 sp61 3183.098862
Rwpos15_62 in15 sp62 11140.846016
Rwpos15_63 in15 sp63 3183.098862
Rwpos15_64 in15 sp64 3183.098862
Rwpos15_65 in15 sp65 3183.098862
Rwpos15_66 in15 sp66 11140.846016
Rwpos15_67 in15 sp67 11140.846016
Rwpos15_68 in15 sp68 3183.098862
Rwpos15_69 in15 sp69 3183.098862
Rwpos15_70 in15 sp70 3183.098862
Rwpos15_71 in15 sp71 3183.098862
Rwpos15_72 in15 sp72 11140.846016
Rwpos15_73 in15 sp73 3183.098862
Rwpos15_74 in15 sp74 11140.846016
Rwpos15_75 in15 sp75 3183.098862
Rwpos15_76 in15 sp76 11140.846016
Rwpos15_77 in15 sp77 11140.846016
Rwpos15_78 in15 sp78 11140.846016
Rwpos15_79 in15 sp79 3183.098862
Rwpos15_80 in15 sp80 3183.098862
Rwpos15_81 in15 sp81 3183.098862
Rwpos15_82 in15 sp82 3183.098862
Rwpos15_83 in15 sp83 3183.098862
Rwpos15_84 in15 sp84 11140.846016
Rwpos15_85 in15 sp85 11140.846016
Rwpos15_86 in15 sp86 11140.846016
Rwpos15_87 in15 sp87 11140.846016
Rwpos15_88 in15 sp88 11140.846016
Rwpos15_89 in15 sp89 3183.098862
Rwpos15_90 in15 sp90 11140.846016
Rwpos15_91 in15 sp91 3183.098862
Rwpos15_92 in15 sp92 3183.098862
Rwpos15_93 in15 sp93 11140.846016
Rwpos15_94 in15 sp94 3183.098862
Rwpos15_95 in15 sp95 3183.098862
Rwpos15_96 in15 sp96 3183.098862
Rwpos15_97 in15 sp97 11140.846016
Rwpos15_98 in15 sp98 3183.098862
Rwpos15_99 in15 sp99 11140.846016
Rwpos15_100 in15 sp100 3183.098862
Rwpos16_1 in16 sp1 3183.098862
Rwpos16_2 in16 sp2 3183.098862
Rwpos16_3 in16 sp3 11140.846016
Rwpos16_4 in16 sp4 11140.846016
Rwpos16_5 in16 sp5 3183.098862
Rwpos16_6 in16 sp6 3183.098862
Rwpos16_7 in16 sp7 11140.846016
Rwpos16_8 in16 sp8 11140.846016
Rwpos16_9 in16 sp9 3183.098862
Rwpos16_10 in16 sp10 11140.846016
Rwpos16_11 in16 sp11 11140.846016
Rwpos16_12 in16 sp12 3183.098862
Rwpos16_13 in16 sp13 3183.098862
Rwpos16_14 in16 sp14 3183.098862
Rwpos16_15 in16 sp15 11140.846016
Rwpos16_16 in16 sp16 3183.098862
Rwpos16_17 in16 sp17 3183.098862
Rwpos16_18 in16 sp18 3183.098862
Rwpos16_19 in16 sp19 11140.846016
Rwpos16_20 in16 sp20 3183.098862
Rwpos16_21 in16 sp21 11140.846016
Rwpos16_22 in16 sp22 3183.098862
Rwpos16_23 in16 sp23 3183.098862
Rwpos16_24 in16 sp24 11140.846016
Rwpos16_25 in16 sp25 11140.846016
Rwpos16_26 in16 sp26 11140.846016
Rwpos16_27 in16 sp27 11140.846016
Rwpos16_28 in16 sp28 11140.846016
Rwpos16_29 in16 sp29 11140.846016
Rwpos16_30 in16 sp30 11140.846016
Rwpos16_31 in16 sp31 11140.846016
Rwpos16_32 in16 sp32 11140.846016
Rwpos16_33 in16 sp33 11140.846016
Rwpos16_34 in16 sp34 11140.846016
Rwpos16_35 in16 sp35 3183.098862
Rwpos16_36 in16 sp36 11140.846016
Rwpos16_37 in16 sp37 11140.846016
Rwpos16_38 in16 sp38 3183.098862
Rwpos16_39 in16 sp39 11140.846016
Rwpos16_40 in16 sp40 3183.098862
Rwpos16_41 in16 sp41 11140.846016
Rwpos16_42 in16 sp42 3183.098862
Rwpos16_43 in16 sp43 11140.846016
Rwpos16_44 in16 sp44 3183.098862
Rwpos16_45 in16 sp45 3183.098862
Rwpos16_46 in16 sp46 11140.846016
Rwpos16_47 in16 sp47 11140.846016
Rwpos16_48 in16 sp48 3183.098862
Rwpos16_49 in16 sp49 3183.098862
Rwpos16_50 in16 sp50 3183.098862
Rwpos16_51 in16 sp51 3183.098862
Rwpos16_52 in16 sp52 11140.846016
Rwpos16_53 in16 sp53 11140.846016
Rwpos16_54 in16 sp54 3183.098862
Rwpos16_55 in16 sp55 11140.846016
Rwpos16_56 in16 sp56 3183.098862
Rwpos16_57 in16 sp57 3183.098862
Rwpos16_58 in16 sp58 11140.846016
Rwpos16_59 in16 sp59 3183.098862
Rwpos16_60 in16 sp60 3183.098862
Rwpos16_61 in16 sp61 3183.098862
Rwpos16_62 in16 sp62 3183.098862
Rwpos16_63 in16 sp63 11140.846016
Rwpos16_64 in16 sp64 11140.846016
Rwpos16_65 in16 sp65 3183.098862
Rwpos16_66 in16 sp66 3183.098862
Rwpos16_67 in16 sp67 3183.098862
Rwpos16_68 in16 sp68 3183.098862
Rwpos16_69 in16 sp69 11140.846016
Rwpos16_70 in16 sp70 3183.098862
Rwpos16_71 in16 sp71 3183.098862
Rwpos16_72 in16 sp72 3183.098862
Rwpos16_73 in16 sp73 3183.098862
Rwpos16_74 in16 sp74 11140.846016
Rwpos16_75 in16 sp75 11140.846016
Rwpos16_76 in16 sp76 3183.098862
Rwpos16_77 in16 sp77 3183.098862
Rwpos16_78 in16 sp78 3183.098862
Rwpos16_79 in16 sp79 11140.846016
Rwpos16_80 in16 sp80 11140.846016
Rwpos16_81 in16 sp81 3183.098862
Rwpos16_82 in16 sp82 3183.098862
Rwpos16_83 in16 sp83 11140.846016
Rwpos16_84 in16 sp84 11140.846016
Rwpos16_85 in16 sp85 11140.846016
Rwpos16_86 in16 sp86 3183.098862
Rwpos16_87 in16 sp87 3183.098862
Rwpos16_88 in16 sp88 3183.098862
Rwpos16_89 in16 sp89 11140.846016
Rwpos16_90 in16 sp90 11140.846016
Rwpos16_91 in16 sp91 11140.846016
Rwpos16_92 in16 sp92 3183.098862
Rwpos16_93 in16 sp93 3183.098862
Rwpos16_94 in16 sp94 11140.846016
Rwpos16_95 in16 sp95 11140.846016
Rwpos16_96 in16 sp96 3183.098862
Rwpos16_97 in16 sp97 3183.098862
Rwpos16_98 in16 sp98 3183.098862
Rwpos16_99 in16 sp99 3183.098862
Rwpos16_100 in16 sp100 11140.846016
Rwpos17_1 in17 sp1 11140.846016
Rwpos17_2 in17 sp2 3183.098862
Rwpos17_3 in17 sp3 11140.846016
Rwpos17_4 in17 sp4 11140.846016
Rwpos17_5 in17 sp5 11140.846016
Rwpos17_6 in17 sp6 11140.846016
Rwpos17_7 in17 sp7 3183.098862
Rwpos17_8 in17 sp8 3183.098862
Rwpos17_9 in17 sp9 3183.098862
Rwpos17_10 in17 sp10 11140.846016
Rwpos17_11 in17 sp11 3183.098862
Rwpos17_12 in17 sp12 3183.098862
Rwpos17_13 in17 sp13 3183.098862
Rwpos17_14 in17 sp14 3183.098862
Rwpos17_15 in17 sp15 3183.098862
Rwpos17_16 in17 sp16 11140.846016
Rwpos17_17 in17 sp17 3183.098862
Rwpos17_18 in17 sp18 3183.098862
Rwpos17_19 in17 sp19 11140.846016
Rwpos17_20 in17 sp20 11140.846016
Rwpos17_21 in17 sp21 11140.846016
Rwpos17_22 in17 sp22 11140.846016
Rwpos17_23 in17 sp23 3183.098862
Rwpos17_24 in17 sp24 3183.098862
Rwpos17_25 in17 sp25 3183.098862
Rwpos17_26 in17 sp26 3183.098862
Rwpos17_27 in17 sp27 11140.846016
Rwpos17_28 in17 sp28 3183.098862
Rwpos17_29 in17 sp29 3183.098862
Rwpos17_30 in17 sp30 3183.098862
Rwpos17_31 in17 sp31 11140.846016
Rwpos17_32 in17 sp32 11140.846016
Rwpos17_33 in17 sp33 3183.098862
Rwpos17_34 in17 sp34 3183.098862
Rwpos17_35 in17 sp35 11140.846016
Rwpos17_36 in17 sp36 3183.098862
Rwpos17_37 in17 sp37 11140.846016
Rwpos17_38 in17 sp38 11140.846016
Rwpos17_39 in17 sp39 3183.098862
Rwpos17_40 in17 sp40 11140.846016
Rwpos17_41 in17 sp41 3183.098862
Rwpos17_42 in17 sp42 11140.846016
Rwpos17_43 in17 sp43 11140.846016
Rwpos17_44 in17 sp44 3183.098862
Rwpos17_45 in17 sp45 3183.098862
Rwpos17_46 in17 sp46 3183.098862
Rwpos17_47 in17 sp47 3183.098862
Rwpos17_48 in17 sp48 11140.846016
Rwpos17_49 in17 sp49 3183.098862
Rwpos17_50 in17 sp50 3183.098862
Rwpos17_51 in17 sp51 11140.846016
Rwpos17_52 in17 sp52 3183.098862
Rwpos17_53 in17 sp53 11140.846016
Rwpos17_54 in17 sp54 11140.846016
Rwpos17_55 in17 sp55 11140.846016
Rwpos17_56 in17 sp56 3183.098862
Rwpos17_57 in17 sp57 3183.098862
Rwpos17_58 in17 sp58 11140.846016
Rwpos17_59 in17 sp59 3183.098862
Rwpos17_60 in17 sp60 3183.098862
Rwpos17_61 in17 sp61 3183.098862
Rwpos17_62 in17 sp62 3183.098862
Rwpos17_63 in17 sp63 3183.098862
Rwpos17_64 in17 sp64 11140.846016
Rwpos17_65 in17 sp65 3183.098862
Rwpos17_66 in17 sp66 11140.846016
Rwpos17_67 in17 sp67 3183.098862
Rwpos17_68 in17 sp68 3183.098862
Rwpos17_69 in17 sp69 11140.846016
Rwpos17_70 in17 sp70 11140.846016
Rwpos17_71 in17 sp71 3183.098862
Rwpos17_72 in17 sp72 3183.098862
Rwpos17_73 in17 sp73 3183.098862
Rwpos17_74 in17 sp74 11140.846016
Rwpos17_75 in17 sp75 3183.098862
Rwpos17_76 in17 sp76 3183.098862
Rwpos17_77 in17 sp77 11140.846016
Rwpos17_78 in17 sp78 3183.098862
Rwpos17_79 in17 sp79 3183.098862
Rwpos17_80 in17 sp80 11140.846016
Rwpos17_81 in17 sp81 11140.846016
Rwpos17_82 in17 sp82 3183.098862
Rwpos17_83 in17 sp83 11140.846016
Rwpos17_84 in17 sp84 3183.098862
Rwpos17_85 in17 sp85 11140.846016
Rwpos17_86 in17 sp86 11140.846016
Rwpos17_87 in17 sp87 3183.098862
Rwpos17_88 in17 sp88 11140.846016
Rwpos17_89 in17 sp89 11140.846016
Rwpos17_90 in17 sp90 11140.846016
Rwpos17_91 in17 sp91 3183.098862
Rwpos17_92 in17 sp92 11140.846016
Rwpos17_93 in17 sp93 3183.098862
Rwpos17_94 in17 sp94 11140.846016
Rwpos17_95 in17 sp95 3183.098862
Rwpos17_96 in17 sp96 11140.846016
Rwpos17_97 in17 sp97 3183.098862
Rwpos17_98 in17 sp98 11140.846016
Rwpos17_99 in17 sp99 11140.846016
Rwpos17_100 in17 sp100 11140.846016
Rwpos18_1 in18 sp1 11140.846016
Rwpos18_2 in18 sp2 11140.846016
Rwpos18_3 in18 sp3 11140.846016
Rwpos18_4 in18 sp4 11140.846016
Rwpos18_5 in18 sp5 11140.846016
Rwpos18_6 in18 sp6 11140.846016
Rwpos18_7 in18 sp7 11140.846016
Rwpos18_8 in18 sp8 3183.098862
Rwpos18_9 in18 sp9 3183.098862
Rwpos18_10 in18 sp10 11140.846016
Rwpos18_11 in18 sp11 11140.846016
Rwpos18_12 in18 sp12 11140.846016
Rwpos18_13 in18 sp13 11140.846016
Rwpos18_14 in18 sp14 11140.846016
Rwpos18_15 in18 sp15 11140.846016
Rwpos18_16 in18 sp16 3183.098862
Rwpos18_17 in18 sp17 3183.098862
Rwpos18_18 in18 sp18 11140.846016
Rwpos18_19 in18 sp19 3183.098862
Rwpos18_20 in18 sp20 11140.846016
Rwpos18_21 in18 sp21 11140.846016
Rwpos18_22 in18 sp22 3183.098862
Rwpos18_23 in18 sp23 3183.098862
Rwpos18_24 in18 sp24 11140.846016
Rwpos18_25 in18 sp25 11140.846016
Rwpos18_26 in18 sp26 3183.098862
Rwpos18_27 in18 sp27 3183.098862
Rwpos18_28 in18 sp28 11140.846016
Rwpos18_29 in18 sp29 3183.098862
Rwpos18_30 in18 sp30 11140.846016
Rwpos18_31 in18 sp31 11140.846016
Rwpos18_32 in18 sp32 11140.846016
Rwpos18_33 in18 sp33 11140.846016
Rwpos18_34 in18 sp34 3183.098862
Rwpos18_35 in18 sp35 3183.098862
Rwpos18_36 in18 sp36 3183.098862
Rwpos18_37 in18 sp37 11140.846016
Rwpos18_38 in18 sp38 3183.098862
Rwpos18_39 in18 sp39 3183.098862
Rwpos18_40 in18 sp40 11140.846016
Rwpos18_41 in18 sp41 11140.846016
Rwpos18_42 in18 sp42 11140.846016
Rwpos18_43 in18 sp43 3183.098862
Rwpos18_44 in18 sp44 11140.846016
Rwpos18_45 in18 sp45 11140.846016
Rwpos18_46 in18 sp46 11140.846016
Rwpos18_47 in18 sp47 3183.098862
Rwpos18_48 in18 sp48 11140.846016
Rwpos18_49 in18 sp49 11140.846016
Rwpos18_50 in18 sp50 11140.846016
Rwpos18_51 in18 sp51 3183.098862
Rwpos18_52 in18 sp52 11140.846016
Rwpos18_53 in18 sp53 3183.098862
Rwpos18_54 in18 sp54 3183.098862
Rwpos18_55 in18 sp55 11140.846016
Rwpos18_56 in18 sp56 3183.098862
Rwpos18_57 in18 sp57 11140.846016
Rwpos18_58 in18 sp58 11140.846016
Rwpos18_59 in18 sp59 11140.846016
Rwpos18_60 in18 sp60 11140.846016
Rwpos18_61 in18 sp61 3183.098862
Rwpos18_62 in18 sp62 3183.098862
Rwpos18_63 in18 sp63 3183.098862
Rwpos18_64 in18 sp64 11140.846016
Rwpos18_65 in18 sp65 3183.098862
Rwpos18_66 in18 sp66 11140.846016
Rwpos18_67 in18 sp67 3183.098862
Rwpos18_68 in18 sp68 11140.846016
Rwpos18_69 in18 sp69 3183.098862
Rwpos18_70 in18 sp70 11140.846016
Rwpos18_71 in18 sp71 11140.846016
Rwpos18_72 in18 sp72 3183.098862
Rwpos18_73 in18 sp73 3183.098862
Rwpos18_74 in18 sp74 11140.846016
Rwpos18_75 in18 sp75 3183.098862
Rwpos18_76 in18 sp76 3183.098862
Rwpos18_77 in18 sp77 3183.098862
Rwpos18_78 in18 sp78 3183.098862
Rwpos18_79 in18 sp79 11140.846016
Rwpos18_80 in18 sp80 3183.098862
Rwpos18_81 in18 sp81 3183.098862
Rwpos18_82 in18 sp82 11140.846016
Rwpos18_83 in18 sp83 11140.846016
Rwpos18_84 in18 sp84 3183.098862
Rwpos18_85 in18 sp85 11140.846016
Rwpos18_86 in18 sp86 11140.846016
Rwpos18_87 in18 sp87 11140.846016
Rwpos18_88 in18 sp88 3183.098862
Rwpos18_89 in18 sp89 11140.846016
Rwpos18_90 in18 sp90 3183.098862
Rwpos18_91 in18 sp91 11140.846016
Rwpos18_92 in18 sp92 11140.846016
Rwpos18_93 in18 sp93 3183.098862
Rwpos18_94 in18 sp94 11140.846016
Rwpos18_95 in18 sp95 11140.846016
Rwpos18_96 in18 sp96 11140.846016
Rwpos18_97 in18 sp97 3183.098862
Rwpos18_98 in18 sp98 3183.098862
Rwpos18_99 in18 sp99 11140.846016
Rwpos18_100 in18 sp100 11140.846016
Rwpos19_1 in19 sp1 3183.098862
Rwpos19_2 in19 sp2 11140.846016
Rwpos19_3 in19 sp3 11140.846016
Rwpos19_4 in19 sp4 11140.846016
Rwpos19_5 in19 sp5 3183.098862
Rwpos19_6 in19 sp6 3183.098862
Rwpos19_7 in19 sp7 11140.846016
Rwpos19_8 in19 sp8 11140.846016
Rwpos19_9 in19 sp9 11140.846016
Rwpos19_10 in19 sp10 3183.098862
Rwpos19_11 in19 sp11 11140.846016
Rwpos19_12 in19 sp12 11140.846016
Rwpos19_13 in19 sp13 3183.098862
Rwpos19_14 in19 sp14 11140.846016
Rwpos19_15 in19 sp15 3183.098862
Rwpos19_16 in19 sp16 3183.098862
Rwpos19_17 in19 sp17 11140.846016
Rwpos19_18 in19 sp18 3183.098862
Rwpos19_19 in19 sp19 11140.846016
Rwpos19_20 in19 sp20 11140.846016
Rwpos19_21 in19 sp21 11140.846016
Rwpos19_22 in19 sp22 11140.846016
Rwpos19_23 in19 sp23 11140.846016
Rwpos19_24 in19 sp24 11140.846016
Rwpos19_25 in19 sp25 3183.098862
Rwpos19_26 in19 sp26 11140.846016
Rwpos19_27 in19 sp27 11140.846016
Rwpos19_28 in19 sp28 11140.846016
Rwpos19_29 in19 sp29 11140.846016
Rwpos19_30 in19 sp30 3183.098862
Rwpos19_31 in19 sp31 11140.846016
Rwpos19_32 in19 sp32 3183.098862
Rwpos19_33 in19 sp33 3183.098862
Rwpos19_34 in19 sp34 3183.098862
Rwpos19_35 in19 sp35 3183.098862
Rwpos19_36 in19 sp36 11140.846016
Rwpos19_37 in19 sp37 11140.846016
Rwpos19_38 in19 sp38 11140.846016
Rwpos19_39 in19 sp39 3183.098862
Rwpos19_40 in19 sp40 11140.846016
Rwpos19_41 in19 sp41 11140.846016
Rwpos19_42 in19 sp42 11140.846016
Rwpos19_43 in19 sp43 11140.846016
Rwpos19_44 in19 sp44 3183.098862
Rwpos19_45 in19 sp45 3183.098862
Rwpos19_46 in19 sp46 3183.098862
Rwpos19_47 in19 sp47 3183.098862
Rwpos19_48 in19 sp48 3183.098862
Rwpos19_49 in19 sp49 3183.098862
Rwpos19_50 in19 sp50 11140.846016
Rwpos19_51 in19 sp51 11140.846016
Rwpos19_52 in19 sp52 3183.098862
Rwpos19_53 in19 sp53 3183.098862
Rwpos19_54 in19 sp54 3183.098862
Rwpos19_55 in19 sp55 3183.098862
Rwpos19_56 in19 sp56 11140.846016
Rwpos19_57 in19 sp57 3183.098862
Rwpos19_58 in19 sp58 11140.846016
Rwpos19_59 in19 sp59 11140.846016
Rwpos19_60 in19 sp60 11140.846016
Rwpos19_61 in19 sp61 3183.098862
Rwpos19_62 in19 sp62 11140.846016
Rwpos19_63 in19 sp63 3183.098862
Rwpos19_64 in19 sp64 3183.098862
Rwpos19_65 in19 sp65 3183.098862
Rwpos19_66 in19 sp66 11140.846016
Rwpos19_67 in19 sp67 11140.846016
Rwpos19_68 in19 sp68 3183.098862
Rwpos19_69 in19 sp69 3183.098862
Rwpos19_70 in19 sp70 11140.846016
Rwpos19_71 in19 sp71 3183.098862
Rwpos19_72 in19 sp72 11140.846016
Rwpos19_73 in19 sp73 11140.846016
Rwpos19_74 in19 sp74 3183.098862
Rwpos19_75 in19 sp75 3183.098862
Rwpos19_76 in19 sp76 3183.098862
Rwpos19_77 in19 sp77 11140.846016
Rwpos19_78 in19 sp78 3183.098862
Rwpos19_79 in19 sp79 3183.098862
Rwpos19_80 in19 sp80 3183.098862
Rwpos19_81 in19 sp81 11140.846016
Rwpos19_82 in19 sp82 3183.098862
Rwpos19_83 in19 sp83 11140.846016
Rwpos19_84 in19 sp84 3183.098862
Rwpos19_85 in19 sp85 3183.098862
Rwpos19_86 in19 sp86 3183.098862
Rwpos19_87 in19 sp87 11140.846016
Rwpos19_88 in19 sp88 11140.846016
Rwpos19_89 in19 sp89 11140.846016
Rwpos19_90 in19 sp90 3183.098862
Rwpos19_91 in19 sp91 11140.846016
Rwpos19_92 in19 sp92 3183.098862
Rwpos19_93 in19 sp93 11140.846016
Rwpos19_94 in19 sp94 3183.098862
Rwpos19_95 in19 sp95 3183.098862
Rwpos19_96 in19 sp96 11140.846016
Rwpos19_97 in19 sp97 11140.846016
Rwpos19_98 in19 sp98 3183.098862
Rwpos19_99 in19 sp99 11140.846016
Rwpos19_100 in19 sp100 11140.846016
Rwpos20_1 in20 sp1 3183.098862
Rwpos20_2 in20 sp2 3183.098862
Rwpos20_3 in20 sp3 11140.846016
Rwpos20_4 in20 sp4 11140.846016
Rwpos20_5 in20 sp5 11140.846016
Rwpos20_6 in20 sp6 11140.846016
Rwpos20_7 in20 sp7 3183.098862
Rwpos20_8 in20 sp8 11140.846016
Rwpos20_9 in20 sp9 11140.846016
Rwpos20_10 in20 sp10 11140.846016
Rwpos20_11 in20 sp11 3183.098862
Rwpos20_12 in20 sp12 11140.846016
Rwpos20_13 in20 sp13 3183.098862
Rwpos20_14 in20 sp14 3183.098862
Rwpos20_15 in20 sp15 11140.846016
Rwpos20_16 in20 sp16 11140.846016
Rwpos20_17 in20 sp17 11140.846016
Rwpos20_18 in20 sp18 3183.098862
Rwpos20_19 in20 sp19 11140.846016
Rwpos20_20 in20 sp20 3183.098862
Rwpos20_21 in20 sp21 11140.846016
Rwpos20_22 in20 sp22 3183.098862
Rwpos20_23 in20 sp23 11140.846016
Rwpos20_24 in20 sp24 3183.098862
Rwpos20_25 in20 sp25 3183.098862
Rwpos20_26 in20 sp26 3183.098862
Rwpos20_27 in20 sp27 3183.098862
Rwpos20_28 in20 sp28 11140.846016
Rwpos20_29 in20 sp29 11140.846016
Rwpos20_30 in20 sp30 11140.846016
Rwpos20_31 in20 sp31 11140.846016
Rwpos20_32 in20 sp32 3183.098862
Rwpos20_33 in20 sp33 3183.098862
Rwpos20_34 in20 sp34 3183.098862
Rwpos20_35 in20 sp35 3183.098862
Rwpos20_36 in20 sp36 11140.846016
Rwpos20_37 in20 sp37 3183.098862
Rwpos20_38 in20 sp38 3183.098862
Rwpos20_39 in20 sp39 11140.846016
Rwpos20_40 in20 sp40 3183.098862
Rwpos20_41 in20 sp41 11140.846016
Rwpos20_42 in20 sp42 11140.846016
Rwpos20_43 in20 sp43 3183.098862
Rwpos20_44 in20 sp44 3183.098862
Rwpos20_45 in20 sp45 3183.098862
Rwpos20_46 in20 sp46 3183.098862
Rwpos20_47 in20 sp47 11140.846016
Rwpos20_48 in20 sp48 3183.098862
Rwpos20_49 in20 sp49 3183.098862
Rwpos20_50 in20 sp50 3183.098862
Rwpos20_51 in20 sp51 3183.098862
Rwpos20_52 in20 sp52 11140.846016
Rwpos20_53 in20 sp53 11140.846016
Rwpos20_54 in20 sp54 3183.098862
Rwpos20_55 in20 sp55 3183.098862
Rwpos20_56 in20 sp56 3183.098862
Rwpos20_57 in20 sp57 11140.846016
Rwpos20_58 in20 sp58 3183.098862
Rwpos20_59 in20 sp59 3183.098862
Rwpos20_60 in20 sp60 11140.846016
Rwpos20_61 in20 sp61 3183.098862
Rwpos20_62 in20 sp62 3183.098862
Rwpos20_63 in20 sp63 11140.846016
Rwpos20_64 in20 sp64 11140.846016
Rwpos20_65 in20 sp65 11140.846016
Rwpos20_66 in20 sp66 3183.098862
Rwpos20_67 in20 sp67 11140.846016
Rwpos20_68 in20 sp68 11140.846016
Rwpos20_69 in20 sp69 11140.846016
Rwpos20_70 in20 sp70 3183.098862
Rwpos20_71 in20 sp71 3183.098862
Rwpos20_72 in20 sp72 3183.098862
Rwpos20_73 in20 sp73 3183.098862
Rwpos20_74 in20 sp74 3183.098862
Rwpos20_75 in20 sp75 3183.098862
Rwpos20_76 in20 sp76 3183.098862
Rwpos20_77 in20 sp77 3183.098862
Rwpos20_78 in20 sp78 3183.098862
Rwpos20_79 in20 sp79 11140.846016
Rwpos20_80 in20 sp80 3183.098862
Rwpos20_81 in20 sp81 3183.098862
Rwpos20_82 in20 sp82 11140.846016
Rwpos20_83 in20 sp83 3183.098862
Rwpos20_84 in20 sp84 3183.098862
Rwpos20_85 in20 sp85 11140.846016
Rwpos20_86 in20 sp86 3183.098862
Rwpos20_87 in20 sp87 3183.098862
Rwpos20_88 in20 sp88 11140.846016
Rwpos20_89 in20 sp89 11140.846016
Rwpos20_90 in20 sp90 3183.098862
Rwpos20_91 in20 sp91 3183.098862
Rwpos20_92 in20 sp92 3183.098862
Rwpos20_93 in20 sp93 3183.098862
Rwpos20_94 in20 sp94 3183.098862
Rwpos20_95 in20 sp95 11140.846016
Rwpos20_96 in20 sp96 11140.846016
Rwpos20_97 in20 sp97 3183.098862
Rwpos20_98 in20 sp98 3183.098862
Rwpos20_99 in20 sp99 3183.098862
Rwpos20_100 in20 sp100 11140.846016
Rwpos21_1 in21 sp1 11140.846016
Rwpos21_2 in21 sp2 3183.098862
Rwpos21_3 in21 sp3 3183.098862
Rwpos21_4 in21 sp4 11140.846016
Rwpos21_5 in21 sp5 3183.098862
Rwpos21_6 in21 sp6 3183.098862
Rwpos21_7 in21 sp7 3183.098862
Rwpos21_8 in21 sp8 3183.098862
Rwpos21_9 in21 sp9 3183.098862
Rwpos21_10 in21 sp10 3183.098862
Rwpos21_11 in21 sp11 11140.846016
Rwpos21_12 in21 sp12 11140.846016
Rwpos21_13 in21 sp13 3183.098862
Rwpos21_14 in21 sp14 11140.846016
Rwpos21_15 in21 sp15 11140.846016
Rwpos21_16 in21 sp16 11140.846016
Rwpos21_17 in21 sp17 3183.098862
Rwpos21_18 in21 sp18 3183.098862
Rwpos21_19 in21 sp19 3183.098862
Rwpos21_20 in21 sp20 11140.846016
Rwpos21_21 in21 sp21 11140.846016
Rwpos21_22 in21 sp22 3183.098862
Rwpos21_23 in21 sp23 3183.098862
Rwpos21_24 in21 sp24 3183.098862
Rwpos21_25 in21 sp25 3183.098862
Rwpos21_26 in21 sp26 3183.098862
Rwpos21_27 in21 sp27 11140.846016
Rwpos21_28 in21 sp28 3183.098862
Rwpos21_29 in21 sp29 3183.098862
Rwpos21_30 in21 sp30 3183.098862
Rwpos21_31 in21 sp31 11140.846016
Rwpos21_32 in21 sp32 11140.846016
Rwpos21_33 in21 sp33 11140.846016
Rwpos21_34 in21 sp34 3183.098862
Rwpos21_35 in21 sp35 3183.098862
Rwpos21_36 in21 sp36 3183.098862
Rwpos21_37 in21 sp37 3183.098862
Rwpos21_38 in21 sp38 3183.098862
Rwpos21_39 in21 sp39 3183.098862
Rwpos21_40 in21 sp40 3183.098862
Rwpos21_41 in21 sp41 11140.846016
Rwpos21_42 in21 sp42 3183.098862
Rwpos21_43 in21 sp43 11140.846016
Rwpos21_44 in21 sp44 3183.098862
Rwpos21_45 in21 sp45 11140.846016
Rwpos21_46 in21 sp46 11140.846016
Rwpos21_47 in21 sp47 11140.846016
Rwpos21_48 in21 sp48 3183.098862
Rwpos21_49 in21 sp49 11140.846016
Rwpos21_50 in21 sp50 3183.098862
Rwpos21_51 in21 sp51 3183.098862
Rwpos21_52 in21 sp52 11140.846016
Rwpos21_53 in21 sp53 11140.846016
Rwpos21_54 in21 sp54 11140.846016
Rwpos21_55 in21 sp55 3183.098862
Rwpos21_56 in21 sp56 3183.098862
Rwpos21_57 in21 sp57 11140.846016
Rwpos21_58 in21 sp58 11140.846016
Rwpos21_59 in21 sp59 11140.846016
Rwpos21_60 in21 sp60 11140.846016
Rwpos21_61 in21 sp61 3183.098862
Rwpos21_62 in21 sp62 3183.098862
Rwpos21_63 in21 sp63 3183.098862
Rwpos21_64 in21 sp64 3183.098862
Rwpos21_65 in21 sp65 11140.846016
Rwpos21_66 in21 sp66 3183.098862
Rwpos21_67 in21 sp67 3183.098862
Rwpos21_68 in21 sp68 3183.098862
Rwpos21_69 in21 sp69 3183.098862
Rwpos21_70 in21 sp70 3183.098862
Rwpos21_71 in21 sp71 11140.846016
Rwpos21_72 in21 sp72 3183.098862
Rwpos21_73 in21 sp73 3183.098862
Rwpos21_74 in21 sp74 3183.098862
Rwpos21_75 in21 sp75 3183.098862
Rwpos21_76 in21 sp76 11140.846016
Rwpos21_77 in21 sp77 3183.098862
Rwpos21_78 in21 sp78 3183.098862
Rwpos21_79 in21 sp79 11140.846016
Rwpos21_80 in21 sp80 11140.846016
Rwpos21_81 in21 sp81 3183.098862
Rwpos21_82 in21 sp82 3183.098862
Rwpos21_83 in21 sp83 3183.098862
Rwpos21_84 in21 sp84 11140.846016
Rwpos21_85 in21 sp85 3183.098862
Rwpos21_86 in21 sp86 11140.846016
Rwpos21_87 in21 sp87 3183.098862
Rwpos21_88 in21 sp88 3183.098862
Rwpos21_89 in21 sp89 3183.098862
Rwpos21_90 in21 sp90 11140.846016
Rwpos21_91 in21 sp91 11140.846016
Rwpos21_92 in21 sp92 3183.098862
Rwpos21_93 in21 sp93 3183.098862
Rwpos21_94 in21 sp94 3183.098862
Rwpos21_95 in21 sp95 3183.098862
Rwpos21_96 in21 sp96 11140.846016
Rwpos21_97 in21 sp97 11140.846016
Rwpos21_98 in21 sp98 3183.098862
Rwpos21_99 in21 sp99 3183.098862
Rwpos21_100 in21 sp100 11140.846016
Rwpos22_1 in22 sp1 3183.098862
Rwpos22_2 in22 sp2 11140.846016
Rwpos22_3 in22 sp3 3183.098862
Rwpos22_4 in22 sp4 3183.098862
Rwpos22_5 in22 sp5 3183.098862
Rwpos22_6 in22 sp6 11140.846016
Rwpos22_7 in22 sp7 11140.846016
Rwpos22_8 in22 sp8 3183.098862
Rwpos22_9 in22 sp9 3183.098862
Rwpos22_10 in22 sp10 3183.098862
Rwpos22_11 in22 sp11 11140.846016
Rwpos22_12 in22 sp12 11140.846016
Rwpos22_13 in22 sp13 11140.846016
Rwpos22_14 in22 sp14 3183.098862
Rwpos22_15 in22 sp15 3183.098862
Rwpos22_16 in22 sp16 11140.846016
Rwpos22_17 in22 sp17 3183.098862
Rwpos22_18 in22 sp18 11140.846016
Rwpos22_19 in22 sp19 3183.098862
Rwpos22_20 in22 sp20 11140.846016
Rwpos22_21 in22 sp21 11140.846016
Rwpos22_22 in22 sp22 11140.846016
Rwpos22_23 in22 sp23 3183.098862
Rwpos22_24 in22 sp24 3183.098862
Rwpos22_25 in22 sp25 3183.098862
Rwpos22_26 in22 sp26 3183.098862
Rwpos22_27 in22 sp27 3183.098862
Rwpos22_28 in22 sp28 11140.846016
Rwpos22_29 in22 sp29 3183.098862
Rwpos22_30 in22 sp30 3183.098862
Rwpos22_31 in22 sp31 11140.846016
Rwpos22_32 in22 sp32 11140.846016
Rwpos22_33 in22 sp33 3183.098862
Rwpos22_34 in22 sp34 11140.846016
Rwpos22_35 in22 sp35 11140.846016
Rwpos22_36 in22 sp36 3183.098862
Rwpos22_37 in22 sp37 3183.098862
Rwpos22_38 in22 sp38 11140.846016
Rwpos22_39 in22 sp39 3183.098862
Rwpos22_40 in22 sp40 3183.098862
Rwpos22_41 in22 sp41 3183.098862
Rwpos22_42 in22 sp42 3183.098862
Rwpos22_43 in22 sp43 11140.846016
Rwpos22_44 in22 sp44 3183.098862
Rwpos22_45 in22 sp45 3183.098862
Rwpos22_46 in22 sp46 11140.846016
Rwpos22_47 in22 sp47 11140.846016
Rwpos22_48 in22 sp48 11140.846016
Rwpos22_49 in22 sp49 11140.846016
Rwpos22_50 in22 sp50 3183.098862
Rwpos22_51 in22 sp51 11140.846016
Rwpos22_52 in22 sp52 11140.846016
Rwpos22_53 in22 sp53 11140.846016
Rwpos22_54 in22 sp54 3183.098862
Rwpos22_55 in22 sp55 11140.846016
Rwpos22_56 in22 sp56 3183.098862
Rwpos22_57 in22 sp57 11140.846016
Rwpos22_58 in22 sp58 3183.098862
Rwpos22_59 in22 sp59 11140.846016
Rwpos22_60 in22 sp60 11140.846016
Rwpos22_61 in22 sp61 11140.846016
Rwpos22_62 in22 sp62 3183.098862
Rwpos22_63 in22 sp63 3183.098862
Rwpos22_64 in22 sp64 11140.846016
Rwpos22_65 in22 sp65 3183.098862
Rwpos22_66 in22 sp66 11140.846016
Rwpos22_67 in22 sp67 11140.846016
Rwpos22_68 in22 sp68 3183.098862
Rwpos22_69 in22 sp69 11140.846016
Rwpos22_70 in22 sp70 11140.846016
Rwpos22_71 in22 sp71 3183.098862
Rwpos22_72 in22 sp72 11140.846016
Rwpos22_73 in22 sp73 11140.846016
Rwpos22_74 in22 sp74 3183.098862
Rwpos22_75 in22 sp75 11140.846016
Rwpos22_76 in22 sp76 11140.846016
Rwpos22_77 in22 sp77 3183.098862
Rwpos22_78 in22 sp78 11140.846016
Rwpos22_79 in22 sp79 11140.846016
Rwpos22_80 in22 sp80 3183.098862
Rwpos22_81 in22 sp81 3183.098862
Rwpos22_82 in22 sp82 3183.098862
Rwpos22_83 in22 sp83 11140.846016
Rwpos22_84 in22 sp84 11140.846016
Rwpos22_85 in22 sp85 11140.846016
Rwpos22_86 in22 sp86 3183.098862
Rwpos22_87 in22 sp87 3183.098862
Rwpos22_88 in22 sp88 3183.098862
Rwpos22_89 in22 sp89 11140.846016
Rwpos22_90 in22 sp90 11140.846016
Rwpos22_91 in22 sp91 3183.098862
Rwpos22_92 in22 sp92 3183.098862
Rwpos22_93 in22 sp93 3183.098862
Rwpos22_94 in22 sp94 11140.846016
Rwpos22_95 in22 sp95 3183.098862
Rwpos22_96 in22 sp96 3183.098862
Rwpos22_97 in22 sp97 3183.098862
Rwpos22_98 in22 sp98 3183.098862
Rwpos22_99 in22 sp99 3183.098862
Rwpos22_100 in22 sp100 3183.098862
Rwpos23_1 in23 sp1 11140.846016
Rwpos23_2 in23 sp2 11140.846016
Rwpos23_3 in23 sp3 11140.846016
Rwpos23_4 in23 sp4 11140.846016
Rwpos23_5 in23 sp5 11140.846016
Rwpos23_6 in23 sp6 3183.098862
Rwpos23_7 in23 sp7 3183.098862
Rwpos23_8 in23 sp8 11140.846016
Rwpos23_9 in23 sp9 11140.846016
Rwpos23_10 in23 sp10 11140.846016
Rwpos23_11 in23 sp11 3183.098862
Rwpos23_12 in23 sp12 3183.098862
Rwpos23_13 in23 sp13 11140.846016
Rwpos23_14 in23 sp14 11140.846016
Rwpos23_15 in23 sp15 3183.098862
Rwpos23_16 in23 sp16 3183.098862
Rwpos23_17 in23 sp17 3183.098862
Rwpos23_18 in23 sp18 11140.846016
Rwpos23_19 in23 sp19 11140.846016
Rwpos23_20 in23 sp20 3183.098862
Rwpos23_21 in23 sp21 3183.098862
Rwpos23_22 in23 sp22 3183.098862
Rwpos23_23 in23 sp23 11140.846016
Rwpos23_24 in23 sp24 11140.846016
Rwpos23_25 in23 sp25 11140.846016
Rwpos23_26 in23 sp26 11140.846016
Rwpos23_27 in23 sp27 3183.098862
Rwpos23_28 in23 sp28 11140.846016
Rwpos23_29 in23 sp29 3183.098862
Rwpos23_30 in23 sp30 3183.098862
Rwpos23_31 in23 sp31 11140.846016
Rwpos23_32 in23 sp32 11140.846016
Rwpos23_33 in23 sp33 3183.098862
Rwpos23_34 in23 sp34 11140.846016
Rwpos23_35 in23 sp35 3183.098862
Rwpos23_36 in23 sp36 3183.098862
Rwpos23_37 in23 sp37 3183.098862
Rwpos23_38 in23 sp38 11140.846016
Rwpos23_39 in23 sp39 11140.846016
Rwpos23_40 in23 sp40 11140.846016
Rwpos23_41 in23 sp41 3183.098862
Rwpos23_42 in23 sp42 11140.846016
Rwpos23_43 in23 sp43 11140.846016
Rwpos23_44 in23 sp44 3183.098862
Rwpos23_45 in23 sp45 11140.846016
Rwpos23_46 in23 sp46 3183.098862
Rwpos23_47 in23 sp47 11140.846016
Rwpos23_48 in23 sp48 11140.846016
Rwpos23_49 in23 sp49 11140.846016
Rwpos23_50 in23 sp50 11140.846016
Rwpos23_51 in23 sp51 3183.098862
Rwpos23_52 in23 sp52 11140.846016
Rwpos23_53 in23 sp53 11140.846016
Rwpos23_54 in23 sp54 3183.098862
Rwpos23_55 in23 sp55 11140.846016
Rwpos23_56 in23 sp56 11140.846016
Rwpos23_57 in23 sp57 11140.846016
Rwpos23_58 in23 sp58 11140.846016
Rwpos23_59 in23 sp59 3183.098862
Rwpos23_60 in23 sp60 3183.098862
Rwpos23_61 in23 sp61 3183.098862
Rwpos23_62 in23 sp62 3183.098862
Rwpos23_63 in23 sp63 11140.846016
Rwpos23_64 in23 sp64 11140.846016
Rwpos23_65 in23 sp65 3183.098862
Rwpos23_66 in23 sp66 3183.098862
Rwpos23_67 in23 sp67 3183.098862
Rwpos23_68 in23 sp68 3183.098862
Rwpos23_69 in23 sp69 11140.846016
Rwpos23_70 in23 sp70 3183.098862
Rwpos23_71 in23 sp71 3183.098862
Rwpos23_72 in23 sp72 11140.846016
Rwpos23_73 in23 sp73 3183.098862
Rwpos23_74 in23 sp74 11140.846016
Rwpos23_75 in23 sp75 11140.846016
Rwpos23_76 in23 sp76 3183.098862
Rwpos23_77 in23 sp77 3183.098862
Rwpos23_78 in23 sp78 3183.098862
Rwpos23_79 in23 sp79 11140.846016
Rwpos23_80 in23 sp80 3183.098862
Rwpos23_81 in23 sp81 11140.846016
Rwpos23_82 in23 sp82 11140.846016
Rwpos23_83 in23 sp83 11140.846016
Rwpos23_84 in23 sp84 11140.846016
Rwpos23_85 in23 sp85 11140.846016
Rwpos23_86 in23 sp86 3183.098862
Rwpos23_87 in23 sp87 11140.846016
Rwpos23_88 in23 sp88 11140.846016
Rwpos23_89 in23 sp89 11140.846016
Rwpos23_90 in23 sp90 3183.098862
Rwpos23_91 in23 sp91 11140.846016
Rwpos23_92 in23 sp92 3183.098862
Rwpos23_93 in23 sp93 11140.846016
Rwpos23_94 in23 sp94 11140.846016
Rwpos23_95 in23 sp95 3183.098862
Rwpos23_96 in23 sp96 11140.846016
Rwpos23_97 in23 sp97 11140.846016
Rwpos23_98 in23 sp98 11140.846016
Rwpos23_99 in23 sp99 3183.098862
Rwpos23_100 in23 sp100 3183.098862
Rwpos24_1 in24 sp1 11140.846016
Rwpos24_2 in24 sp2 3183.098862
Rwpos24_3 in24 sp3 11140.846016
Rwpos24_4 in24 sp4 11140.846016
Rwpos24_5 in24 sp5 11140.846016
Rwpos24_6 in24 sp6 11140.846016
Rwpos24_7 in24 sp7 3183.098862
Rwpos24_8 in24 sp8 11140.846016
Rwpos24_9 in24 sp9 11140.846016
Rwpos24_10 in24 sp10 3183.098862
Rwpos24_11 in24 sp11 11140.846016
Rwpos24_12 in24 sp12 11140.846016
Rwpos24_13 in24 sp13 11140.846016
Rwpos24_14 in24 sp14 11140.846016
Rwpos24_15 in24 sp15 3183.098862
Rwpos24_16 in24 sp16 11140.846016
Rwpos24_17 in24 sp17 11140.846016
Rwpos24_18 in24 sp18 3183.098862
Rwpos24_19 in24 sp19 3183.098862
Rwpos24_20 in24 sp20 11140.846016
Rwpos24_21 in24 sp21 3183.098862
Rwpos24_22 in24 sp22 11140.846016
Rwpos24_23 in24 sp23 11140.846016
Rwpos24_24 in24 sp24 3183.098862
Rwpos24_25 in24 sp25 11140.846016
Rwpos24_26 in24 sp26 3183.098862
Rwpos24_27 in24 sp27 3183.098862
Rwpos24_28 in24 sp28 11140.846016
Rwpos24_29 in24 sp29 11140.846016
Rwpos24_30 in24 sp30 11140.846016
Rwpos24_31 in24 sp31 11140.846016
Rwpos24_32 in24 sp32 3183.098862
Rwpos24_33 in24 sp33 3183.098862
Rwpos24_34 in24 sp34 11140.846016
Rwpos24_35 in24 sp35 3183.098862
Rwpos24_36 in24 sp36 11140.846016
Rwpos24_37 in24 sp37 3183.098862
Rwpos24_38 in24 sp38 11140.846016
Rwpos24_39 in24 sp39 11140.846016
Rwpos24_40 in24 sp40 3183.098862
Rwpos24_41 in24 sp41 11140.846016
Rwpos24_42 in24 sp42 11140.846016
Rwpos24_43 in24 sp43 3183.098862
Rwpos24_44 in24 sp44 11140.846016
Rwpos24_45 in24 sp45 3183.098862
Rwpos24_46 in24 sp46 3183.098862
Rwpos24_47 in24 sp47 11140.846016
Rwpos24_48 in24 sp48 11140.846016
Rwpos24_49 in24 sp49 11140.846016
Rwpos24_50 in24 sp50 11140.846016
Rwpos24_51 in24 sp51 3183.098862
Rwpos24_52 in24 sp52 3183.098862
Rwpos24_53 in24 sp53 11140.846016
Rwpos24_54 in24 sp54 3183.098862
Rwpos24_55 in24 sp55 3183.098862
Rwpos24_56 in24 sp56 3183.098862
Rwpos24_57 in24 sp57 11140.846016
Rwpos24_58 in24 sp58 3183.098862
Rwpos24_59 in24 sp59 11140.846016
Rwpos24_60 in24 sp60 3183.098862
Rwpos24_61 in24 sp61 3183.098862
Rwpos24_62 in24 sp62 3183.098862
Rwpos24_63 in24 sp63 11140.846016
Rwpos24_64 in24 sp64 11140.846016
Rwpos24_65 in24 sp65 11140.846016
Rwpos24_66 in24 sp66 3183.098862
Rwpos24_67 in24 sp67 3183.098862
Rwpos24_68 in24 sp68 3183.098862
Rwpos24_69 in24 sp69 11140.846016
Rwpos24_70 in24 sp70 3183.098862
Rwpos24_71 in24 sp71 3183.098862
Rwpos24_72 in24 sp72 11140.846016
Rwpos24_73 in24 sp73 11140.846016
Rwpos24_74 in24 sp74 11140.846016
Rwpos24_75 in24 sp75 3183.098862
Rwpos24_76 in24 sp76 11140.846016
Rwpos24_77 in24 sp77 3183.098862
Rwpos24_78 in24 sp78 3183.098862
Rwpos24_79 in24 sp79 11140.846016
Rwpos24_80 in24 sp80 3183.098862
Rwpos24_81 in24 sp81 3183.098862
Rwpos24_82 in24 sp82 3183.098862
Rwpos24_83 in24 sp83 3183.098862
Rwpos24_84 in24 sp84 11140.846016
Rwpos24_85 in24 sp85 11140.846016
Rwpos24_86 in24 sp86 3183.098862
Rwpos24_87 in24 sp87 3183.098862
Rwpos24_88 in24 sp88 3183.098862
Rwpos24_89 in24 sp89 3183.098862
Rwpos24_90 in24 sp90 11140.846016
Rwpos24_91 in24 sp91 11140.846016
Rwpos24_92 in24 sp92 3183.098862
Rwpos24_93 in24 sp93 3183.098862
Rwpos24_94 in24 sp94 11140.846016
Rwpos24_95 in24 sp95 11140.846016
Rwpos24_96 in24 sp96 11140.846016
Rwpos24_97 in24 sp97 3183.098862
Rwpos24_98 in24 sp98 3183.098862
Rwpos24_99 in24 sp99 3183.098862
Rwpos24_100 in24 sp100 3183.098862
Rwpos25_1 in25 sp1 3183.098862
Rwpos25_2 in25 sp2 3183.098862
Rwpos25_3 in25 sp3 3183.098862
Rwpos25_4 in25 sp4 3183.098862
Rwpos25_5 in25 sp5 3183.098862
Rwpos25_6 in25 sp6 11140.846016
Rwpos25_7 in25 sp7 3183.098862
Rwpos25_8 in25 sp8 11140.846016
Rwpos25_9 in25 sp9 11140.846016
Rwpos25_10 in25 sp10 3183.098862
Rwpos25_11 in25 sp11 11140.846016
Rwpos25_12 in25 sp12 11140.846016
Rwpos25_13 in25 sp13 3183.098862
Rwpos25_14 in25 sp14 11140.846016
Rwpos25_15 in25 sp15 3183.098862
Rwpos25_16 in25 sp16 11140.846016
Rwpos25_17 in25 sp17 11140.846016
Rwpos25_18 in25 sp18 3183.098862
Rwpos25_19 in25 sp19 3183.098862
Rwpos25_20 in25 sp20 3183.098862
Rwpos25_21 in25 sp21 11140.846016
Rwpos25_22 in25 sp22 3183.098862
Rwpos25_23 in25 sp23 3183.098862
Rwpos25_24 in25 sp24 11140.846016
Rwpos25_25 in25 sp25 3183.098862
Rwpos25_26 in25 sp26 3183.098862
Rwpos25_27 in25 sp27 11140.846016
Rwpos25_28 in25 sp28 11140.846016
Rwpos25_29 in25 sp29 3183.098862
Rwpos25_30 in25 sp30 3183.098862
Rwpos25_31 in25 sp31 3183.098862
Rwpos25_32 in25 sp32 11140.846016
Rwpos25_33 in25 sp33 3183.098862
Rwpos25_34 in25 sp34 11140.846016
Rwpos25_35 in25 sp35 3183.098862
Rwpos25_36 in25 sp36 3183.098862
Rwpos25_37 in25 sp37 3183.098862
Rwpos25_38 in25 sp38 11140.846016
Rwpos25_39 in25 sp39 3183.098862
Rwpos25_40 in25 sp40 3183.098862
Rwpos25_41 in25 sp41 3183.098862
Rwpos25_42 in25 sp42 11140.846016
Rwpos25_43 in25 sp43 11140.846016
Rwpos25_44 in25 sp44 3183.098862
Rwpos25_45 in25 sp45 11140.846016
Rwpos25_46 in25 sp46 11140.846016
Rwpos25_47 in25 sp47 3183.098862
Rwpos25_48 in25 sp48 3183.098862
Rwpos25_49 in25 sp49 11140.846016
Rwpos25_50 in25 sp50 11140.846016
Rwpos25_51 in25 sp51 3183.098862
Rwpos25_52 in25 sp52 3183.098862
Rwpos25_53 in25 sp53 3183.098862
Rwpos25_54 in25 sp54 3183.098862
Rwpos25_55 in25 sp55 3183.098862
Rwpos25_56 in25 sp56 3183.098862
Rwpos25_57 in25 sp57 11140.846016
Rwpos25_58 in25 sp58 3183.098862
Rwpos25_59 in25 sp59 11140.846016
Rwpos25_60 in25 sp60 11140.846016
Rwpos25_61 in25 sp61 3183.098862
Rwpos25_62 in25 sp62 3183.098862
Rwpos25_63 in25 sp63 3183.098862
Rwpos25_64 in25 sp64 3183.098862
Rwpos25_65 in25 sp65 3183.098862
Rwpos25_66 in25 sp66 11140.846016
Rwpos25_67 in25 sp67 3183.098862
Rwpos25_68 in25 sp68 3183.098862
Rwpos25_69 in25 sp69 3183.098862
Rwpos25_70 in25 sp70 3183.098862
Rwpos25_71 in25 sp71 3183.098862
Rwpos25_72 in25 sp72 3183.098862
Rwpos25_73 in25 sp73 3183.098862
Rwpos25_74 in25 sp74 3183.098862
Rwpos25_75 in25 sp75 11140.846016
Rwpos25_76 in25 sp76 11140.846016
Rwpos25_77 in25 sp77 11140.846016
Rwpos25_78 in25 sp78 11140.846016
Rwpos25_79 in25 sp79 11140.846016
Rwpos25_80 in25 sp80 3183.098862
Rwpos25_81 in25 sp81 3183.098862
Rwpos25_82 in25 sp82 11140.846016
Rwpos25_83 in25 sp83 3183.098862
Rwpos25_84 in25 sp84 3183.098862
Rwpos25_85 in25 sp85 11140.846016
Rwpos25_86 in25 sp86 11140.846016
Rwpos25_87 in25 sp87 3183.098862
Rwpos25_88 in25 sp88 3183.098862
Rwpos25_89 in25 sp89 3183.098862
Rwpos25_90 in25 sp90 3183.098862
Rwpos25_91 in25 sp91 11140.846016
Rwpos25_92 in25 sp92 11140.846016
Rwpos25_93 in25 sp93 3183.098862
Rwpos25_94 in25 sp94 11140.846016
Rwpos25_95 in25 sp95 11140.846016
Rwpos25_96 in25 sp96 11140.846016
Rwpos25_97 in25 sp97 3183.098862
Rwpos25_98 in25 sp98 11140.846016
Rwpos25_99 in25 sp99 3183.098862
Rwpos25_100 in25 sp100 3183.098862
Rwpos26_1 in26 sp1 3183.098862
Rwpos26_2 in26 sp2 11140.846016
Rwpos26_3 in26 sp3 3183.098862
Rwpos26_4 in26 sp4 3183.098862
Rwpos26_5 in26 sp5 11140.846016
Rwpos26_6 in26 sp6 3183.098862
Rwpos26_7 in26 sp7 11140.846016
Rwpos26_8 in26 sp8 11140.846016
Rwpos26_9 in26 sp9 11140.846016
Rwpos26_10 in26 sp10 11140.846016
Rwpos26_11 in26 sp11 3183.098862
Rwpos26_12 in26 sp12 11140.846016
Rwpos26_13 in26 sp13 3183.098862
Rwpos26_14 in26 sp14 11140.846016
Rwpos26_15 in26 sp15 3183.098862
Rwpos26_16 in26 sp16 3183.098862
Rwpos26_17 in26 sp17 3183.098862
Rwpos26_18 in26 sp18 3183.098862
Rwpos26_19 in26 sp19 3183.098862
Rwpos26_20 in26 sp20 3183.098862
Rwpos26_21 in26 sp21 11140.846016
Rwpos26_22 in26 sp22 3183.098862
Rwpos26_23 in26 sp23 3183.098862
Rwpos26_24 in26 sp24 11140.846016
Rwpos26_25 in26 sp25 11140.846016
Rwpos26_26 in26 sp26 11140.846016
Rwpos26_27 in26 sp27 3183.098862
Rwpos26_28 in26 sp28 3183.098862
Rwpos26_29 in26 sp29 3183.098862
Rwpos26_30 in26 sp30 11140.846016
Rwpos26_31 in26 sp31 3183.098862
Rwpos26_32 in26 sp32 3183.098862
Rwpos26_33 in26 sp33 3183.098862
Rwpos26_34 in26 sp34 11140.846016
Rwpos26_35 in26 sp35 3183.098862
Rwpos26_36 in26 sp36 3183.098862
Rwpos26_37 in26 sp37 11140.846016
Rwpos26_38 in26 sp38 11140.846016
Rwpos26_39 in26 sp39 11140.846016
Rwpos26_40 in26 sp40 11140.846016
Rwpos26_41 in26 sp41 3183.098862
Rwpos26_42 in26 sp42 11140.846016
Rwpos26_43 in26 sp43 11140.846016
Rwpos26_44 in26 sp44 11140.846016
Rwpos26_45 in26 sp45 3183.098862
Rwpos26_46 in26 sp46 3183.098862
Rwpos26_47 in26 sp47 3183.098862
Rwpos26_48 in26 sp48 11140.846016
Rwpos26_49 in26 sp49 3183.098862
Rwpos26_50 in26 sp50 3183.098862
Rwpos26_51 in26 sp51 3183.098862
Rwpos26_52 in26 sp52 3183.098862
Rwpos26_53 in26 sp53 11140.846016
Rwpos26_54 in26 sp54 3183.098862
Rwpos26_55 in26 sp55 3183.098862
Rwpos26_56 in26 sp56 11140.846016
Rwpos26_57 in26 sp57 11140.846016
Rwpos26_58 in26 sp58 3183.098862
Rwpos26_59 in26 sp59 11140.846016
Rwpos26_60 in26 sp60 3183.098862
Rwpos26_61 in26 sp61 3183.098862
Rwpos26_62 in26 sp62 11140.846016
Rwpos26_63 in26 sp63 3183.098862
Rwpos26_64 in26 sp64 11140.846016
Rwpos26_65 in26 sp65 3183.098862
Rwpos26_66 in26 sp66 11140.846016
Rwpos26_67 in26 sp67 11140.846016
Rwpos26_68 in26 sp68 11140.846016
Rwpos26_69 in26 sp69 3183.098862
Rwpos26_70 in26 sp70 11140.846016
Rwpos26_71 in26 sp71 3183.098862
Rwpos26_72 in26 sp72 3183.098862
Rwpos26_73 in26 sp73 11140.846016
Rwpos26_74 in26 sp74 3183.098862
Rwpos26_75 in26 sp75 3183.098862
Rwpos26_76 in26 sp76 11140.846016
Rwpos26_77 in26 sp77 3183.098862
Rwpos26_78 in26 sp78 3183.098862
Rwpos26_79 in26 sp79 3183.098862
Rwpos26_80 in26 sp80 11140.846016
Rwpos26_81 in26 sp81 3183.098862
Rwpos26_82 in26 sp82 3183.098862
Rwpos26_83 in26 sp83 11140.846016
Rwpos26_84 in26 sp84 3183.098862
Rwpos26_85 in26 sp85 11140.846016
Rwpos26_86 in26 sp86 3183.098862
Rwpos26_87 in26 sp87 3183.098862
Rwpos26_88 in26 sp88 11140.846016
Rwpos26_89 in26 sp89 3183.098862
Rwpos26_90 in26 sp90 11140.846016
Rwpos26_91 in26 sp91 11140.846016
Rwpos26_92 in26 sp92 3183.098862
Rwpos26_93 in26 sp93 3183.098862
Rwpos26_94 in26 sp94 11140.846016
Rwpos26_95 in26 sp95 3183.098862
Rwpos26_96 in26 sp96 11140.846016
Rwpos26_97 in26 sp97 3183.098862
Rwpos26_98 in26 sp98 11140.846016
Rwpos26_99 in26 sp99 11140.846016
Rwpos26_100 in26 sp100 3183.098862
Rwpos27_1 in27 sp1 3183.098862
Rwpos27_2 in27 sp2 11140.846016
Rwpos27_3 in27 sp3 3183.098862
Rwpos27_4 in27 sp4 3183.098862
Rwpos27_5 in27 sp5 11140.846016
Rwpos27_6 in27 sp6 3183.098862
Rwpos27_7 in27 sp7 3183.098862
Rwpos27_8 in27 sp8 11140.846016
Rwpos27_9 in27 sp9 3183.098862
Rwpos27_10 in27 sp10 11140.846016
Rwpos27_11 in27 sp11 11140.846016
Rwpos27_12 in27 sp12 11140.846016
Rwpos27_13 in27 sp13 11140.846016
Rwpos27_14 in27 sp14 3183.098862
Rwpos27_15 in27 sp15 11140.846016
Rwpos27_16 in27 sp16 11140.846016
Rwpos27_17 in27 sp17 3183.098862
Rwpos27_18 in27 sp18 11140.846016
Rwpos27_19 in27 sp19 3183.098862
Rwpos27_20 in27 sp20 3183.098862
Rwpos27_21 in27 sp21 11140.846016
Rwpos27_22 in27 sp22 3183.098862
Rwpos27_23 in27 sp23 3183.098862
Rwpos27_24 in27 sp24 11140.846016
Rwpos27_25 in27 sp25 3183.098862
Rwpos27_26 in27 sp26 3183.098862
Rwpos27_27 in27 sp27 3183.098862
Rwpos27_28 in27 sp28 3183.098862
Rwpos27_29 in27 sp29 11140.846016
Rwpos27_30 in27 sp30 3183.098862
Rwpos27_31 in27 sp31 11140.846016
Rwpos27_32 in27 sp32 11140.846016
Rwpos27_33 in27 sp33 11140.846016
Rwpos27_34 in27 sp34 11140.846016
Rwpos27_35 in27 sp35 3183.098862
Rwpos27_36 in27 sp36 3183.098862
Rwpos27_37 in27 sp37 11140.846016
Rwpos27_38 in27 sp38 3183.098862
Rwpos27_39 in27 sp39 3183.098862
Rwpos27_40 in27 sp40 3183.098862
Rwpos27_41 in27 sp41 11140.846016
Rwpos27_42 in27 sp42 3183.098862
Rwpos27_43 in27 sp43 11140.846016
Rwpos27_44 in27 sp44 3183.098862
Rwpos27_45 in27 sp45 3183.098862
Rwpos27_46 in27 sp46 3183.098862
Rwpos27_47 in27 sp47 3183.098862
Rwpos27_48 in27 sp48 3183.098862
Rwpos27_49 in27 sp49 11140.846016
Rwpos27_50 in27 sp50 3183.098862
Rwpos27_51 in27 sp51 3183.098862
Rwpos27_52 in27 sp52 3183.098862
Rwpos27_53 in27 sp53 3183.098862
Rwpos27_54 in27 sp54 11140.846016
Rwpos27_55 in27 sp55 11140.846016
Rwpos27_56 in27 sp56 3183.098862
Rwpos27_57 in27 sp57 11140.846016
Rwpos27_58 in27 sp58 11140.846016
Rwpos27_59 in27 sp59 11140.846016
Rwpos27_60 in27 sp60 11140.846016
Rwpos27_61 in27 sp61 3183.098862
Rwpos27_62 in27 sp62 3183.098862
Rwpos27_63 in27 sp63 3183.098862
Rwpos27_64 in27 sp64 3183.098862
Rwpos27_65 in27 sp65 3183.098862
Rwpos27_66 in27 sp66 11140.846016
Rwpos27_67 in27 sp67 3183.098862
Rwpos27_68 in27 sp68 3183.098862
Rwpos27_69 in27 sp69 3183.098862
Rwpos27_70 in27 sp70 3183.098862
Rwpos27_71 in27 sp71 3183.098862
Rwpos27_72 in27 sp72 3183.098862
Rwpos27_73 in27 sp73 11140.846016
Rwpos27_74 in27 sp74 3183.098862
Rwpos27_75 in27 sp75 11140.846016
Rwpos27_76 in27 sp76 3183.098862
Rwpos27_77 in27 sp77 11140.846016
Rwpos27_78 in27 sp78 3183.098862
Rwpos27_79 in27 sp79 11140.846016
Rwpos27_80 in27 sp80 3183.098862
Rwpos27_81 in27 sp81 3183.098862
Rwpos27_82 in27 sp82 11140.846016
Rwpos27_83 in27 sp83 3183.098862
Rwpos27_84 in27 sp84 11140.846016
Rwpos27_85 in27 sp85 3183.098862
Rwpos27_86 in27 sp86 3183.098862
Rwpos27_87 in27 sp87 11140.846016
Rwpos27_88 in27 sp88 11140.846016
Rwpos27_89 in27 sp89 3183.098862
Rwpos27_90 in27 sp90 3183.098862
Rwpos27_91 in27 sp91 11140.846016
Rwpos27_92 in27 sp92 11140.846016
Rwpos27_93 in27 sp93 11140.846016
Rwpos27_94 in27 sp94 11140.846016
Rwpos27_95 in27 sp95 3183.098862
Rwpos27_96 in27 sp96 3183.098862
Rwpos27_97 in27 sp97 11140.846016
Rwpos27_98 in27 sp98 3183.098862
Rwpos27_99 in27 sp99 3183.098862
Rwpos27_100 in27 sp100 11140.846016
Rwpos28_1 in28 sp1 11140.846016
Rwpos28_2 in28 sp2 11140.846016
Rwpos28_3 in28 sp3 3183.098862
Rwpos28_4 in28 sp4 3183.098862
Rwpos28_5 in28 sp5 3183.098862
Rwpos28_6 in28 sp6 11140.846016
Rwpos28_7 in28 sp7 11140.846016
Rwpos28_8 in28 sp8 3183.098862
Rwpos28_9 in28 sp9 11140.846016
Rwpos28_10 in28 sp10 11140.846016
Rwpos28_11 in28 sp11 11140.846016
Rwpos28_12 in28 sp12 11140.846016
Rwpos28_13 in28 sp13 11140.846016
Rwpos28_14 in28 sp14 3183.098862
Rwpos28_15 in28 sp15 11140.846016
Rwpos28_16 in28 sp16 11140.846016
Rwpos28_17 in28 sp17 3183.098862
Rwpos28_18 in28 sp18 3183.098862
Rwpos28_19 in28 sp19 3183.098862
Rwpos28_20 in28 sp20 11140.846016
Rwpos28_21 in28 sp21 11140.846016
Rwpos28_22 in28 sp22 11140.846016
Rwpos28_23 in28 sp23 11140.846016
Rwpos28_24 in28 sp24 11140.846016
Rwpos28_25 in28 sp25 3183.098862
Rwpos28_26 in28 sp26 3183.098862
Rwpos28_27 in28 sp27 3183.098862
Rwpos28_28 in28 sp28 3183.098862
Rwpos28_29 in28 sp29 11140.846016
Rwpos28_30 in28 sp30 3183.098862
Rwpos28_31 in28 sp31 3183.098862
Rwpos28_32 in28 sp32 3183.098862
Rwpos28_33 in28 sp33 11140.846016
Rwpos28_34 in28 sp34 3183.098862
Rwpos28_35 in28 sp35 3183.098862
Rwpos28_36 in28 sp36 3183.098862
Rwpos28_37 in28 sp37 3183.098862
Rwpos28_38 in28 sp38 11140.846016
Rwpos28_39 in28 sp39 3183.098862
Rwpos28_40 in28 sp40 11140.846016
Rwpos28_41 in28 sp41 3183.098862
Rwpos28_42 in28 sp42 3183.098862
Rwpos28_43 in28 sp43 3183.098862
Rwpos28_44 in28 sp44 11140.846016
Rwpos28_45 in28 sp45 11140.846016
Rwpos28_46 in28 sp46 3183.098862
Rwpos28_47 in28 sp47 11140.846016
Rwpos28_48 in28 sp48 3183.098862
Rwpos28_49 in28 sp49 3183.098862
Rwpos28_50 in28 sp50 3183.098862
Rwpos28_51 in28 sp51 11140.846016
Rwpos28_52 in28 sp52 3183.098862
Rwpos28_53 in28 sp53 3183.098862
Rwpos28_54 in28 sp54 11140.846016
Rwpos28_55 in28 sp55 11140.846016
Rwpos28_56 in28 sp56 11140.846016
Rwpos28_57 in28 sp57 3183.098862
Rwpos28_58 in28 sp58 11140.846016
Rwpos28_59 in28 sp59 11140.846016
Rwpos28_60 in28 sp60 3183.098862
Rwpos28_61 in28 sp61 3183.098862
Rwpos28_62 in28 sp62 3183.098862
Rwpos28_63 in28 sp63 11140.846016
Rwpos28_64 in28 sp64 3183.098862
Rwpos28_65 in28 sp65 3183.098862
Rwpos28_66 in28 sp66 11140.846016
Rwpos28_67 in28 sp67 3183.098862
Rwpos28_68 in28 sp68 3183.098862
Rwpos28_69 in28 sp69 11140.846016
Rwpos28_70 in28 sp70 3183.098862
Rwpos28_71 in28 sp71 11140.846016
Rwpos28_72 in28 sp72 3183.098862
Rwpos28_73 in28 sp73 11140.846016
Rwpos28_74 in28 sp74 11140.846016
Rwpos28_75 in28 sp75 11140.846016
Rwpos28_76 in28 sp76 3183.098862
Rwpos28_77 in28 sp77 3183.098862
Rwpos28_78 in28 sp78 3183.098862
Rwpos28_79 in28 sp79 11140.846016
Rwpos28_80 in28 sp80 3183.098862
Rwpos28_81 in28 sp81 3183.098862
Rwpos28_82 in28 sp82 3183.098862
Rwpos28_83 in28 sp83 3183.098862
Rwpos28_84 in28 sp84 3183.098862
Rwpos28_85 in28 sp85 11140.846016
Rwpos28_86 in28 sp86 11140.846016
Rwpos28_87 in28 sp87 3183.098862
Rwpos28_88 in28 sp88 11140.846016
Rwpos28_89 in28 sp89 3183.098862
Rwpos28_90 in28 sp90 11140.846016
Rwpos28_91 in28 sp91 11140.846016
Rwpos28_92 in28 sp92 11140.846016
Rwpos28_93 in28 sp93 3183.098862
Rwpos28_94 in28 sp94 11140.846016
Rwpos28_95 in28 sp95 11140.846016
Rwpos28_96 in28 sp96 3183.098862
Rwpos28_97 in28 sp97 3183.098862
Rwpos28_98 in28 sp98 3183.098862
Rwpos28_99 in28 sp99 11140.846016
Rwpos28_100 in28 sp100 11140.846016
Rwpos29_1 in29 sp1 3183.098862
Rwpos29_2 in29 sp2 3183.098862
Rwpos29_3 in29 sp3 3183.098862
Rwpos29_4 in29 sp4 11140.846016
Rwpos29_5 in29 sp5 11140.846016
Rwpos29_6 in29 sp6 11140.846016
Rwpos29_7 in29 sp7 3183.098862
Rwpos29_8 in29 sp8 3183.098862
Rwpos29_9 in29 sp9 3183.098862
Rwpos29_10 in29 sp10 11140.846016
Rwpos29_11 in29 sp11 11140.846016
Rwpos29_12 in29 sp12 11140.846016
Rwpos29_13 in29 sp13 3183.098862
Rwpos29_14 in29 sp14 3183.098862
Rwpos29_15 in29 sp15 3183.098862
Rwpos29_16 in29 sp16 11140.846016
Rwpos29_17 in29 sp17 11140.846016
Rwpos29_18 in29 sp18 11140.846016
Rwpos29_19 in29 sp19 3183.098862
Rwpos29_20 in29 sp20 3183.098862
Rwpos29_21 in29 sp21 3183.098862
Rwpos29_22 in29 sp22 3183.098862
Rwpos29_23 in29 sp23 3183.098862
Rwpos29_24 in29 sp24 3183.098862
Rwpos29_25 in29 sp25 3183.098862
Rwpos29_26 in29 sp26 3183.098862
Rwpos29_27 in29 sp27 11140.846016
Rwpos29_28 in29 sp28 3183.098862
Rwpos29_29 in29 sp29 11140.846016
Rwpos29_30 in29 sp30 11140.846016
Rwpos29_31 in29 sp31 11140.846016
Rwpos29_32 in29 sp32 11140.846016
Rwpos29_33 in29 sp33 11140.846016
Rwpos29_34 in29 sp34 3183.098862
Rwpos29_35 in29 sp35 3183.098862
Rwpos29_36 in29 sp36 11140.846016
Rwpos29_37 in29 sp37 11140.846016
Rwpos29_38 in29 sp38 11140.846016
Rwpos29_39 in29 sp39 3183.098862
Rwpos29_40 in29 sp40 3183.098862
Rwpos29_41 in29 sp41 3183.098862
Rwpos29_42 in29 sp42 11140.846016
Rwpos29_43 in29 sp43 11140.846016
Rwpos29_44 in29 sp44 3183.098862
Rwpos29_45 in29 sp45 3183.098862
Rwpos29_46 in29 sp46 3183.098862
Rwpos29_47 in29 sp47 3183.098862
Rwpos29_48 in29 sp48 11140.846016
Rwpos29_49 in29 sp49 11140.846016
Rwpos29_50 in29 sp50 3183.098862
Rwpos29_51 in29 sp51 3183.098862
Rwpos29_52 in29 sp52 3183.098862
Rwpos29_53 in29 sp53 11140.846016
Rwpos29_54 in29 sp54 11140.846016
Rwpos29_55 in29 sp55 3183.098862
Rwpos29_56 in29 sp56 3183.098862
Rwpos29_57 in29 sp57 3183.098862
Rwpos29_58 in29 sp58 3183.098862
Rwpos29_59 in29 sp59 11140.846016
Rwpos29_60 in29 sp60 3183.098862
Rwpos29_61 in29 sp61 11140.846016
Rwpos29_62 in29 sp62 3183.098862
Rwpos29_63 in29 sp63 3183.098862
Rwpos29_64 in29 sp64 3183.098862
Rwpos29_65 in29 sp65 11140.846016
Rwpos29_66 in29 sp66 11140.846016
Rwpos29_67 in29 sp67 3183.098862
Rwpos29_68 in29 sp68 11140.846016
Rwpos29_69 in29 sp69 11140.846016
Rwpos29_70 in29 sp70 11140.846016
Rwpos29_71 in29 sp71 3183.098862
Rwpos29_72 in29 sp72 3183.098862
Rwpos29_73 in29 sp73 3183.098862
Rwpos29_74 in29 sp74 3183.098862
Rwpos29_75 in29 sp75 11140.846016
Rwpos29_76 in29 sp76 11140.846016
Rwpos29_77 in29 sp77 3183.098862
Rwpos29_78 in29 sp78 11140.846016
Rwpos29_79 in29 sp79 11140.846016
Rwpos29_80 in29 sp80 3183.098862
Rwpos29_81 in29 sp81 11140.846016
Rwpos29_82 in29 sp82 11140.846016
Rwpos29_83 in29 sp83 11140.846016
Rwpos29_84 in29 sp84 11140.846016
Rwpos29_85 in29 sp85 3183.098862
Rwpos29_86 in29 sp86 11140.846016
Rwpos29_87 in29 sp87 3183.098862
Rwpos29_88 in29 sp88 3183.098862
Rwpos29_89 in29 sp89 3183.098862
Rwpos29_90 in29 sp90 3183.098862
Rwpos29_91 in29 sp91 11140.846016
Rwpos29_92 in29 sp92 11140.846016
Rwpos29_93 in29 sp93 3183.098862
Rwpos29_94 in29 sp94 3183.098862
Rwpos29_95 in29 sp95 3183.098862
Rwpos29_96 in29 sp96 11140.846016
Rwpos29_97 in29 sp97 3183.098862
Rwpos29_98 in29 sp98 3183.098862
Rwpos29_99 in29 sp99 11140.846016
Rwpos29_100 in29 sp100 3183.098862
Rwpos30_1 in30 sp1 11140.846016
Rwpos30_2 in30 sp2 11140.846016
Rwpos30_3 in30 sp3 3183.098862
Rwpos30_4 in30 sp4 3183.098862
Rwpos30_5 in30 sp5 3183.098862
Rwpos30_6 in30 sp6 3183.098862
Rwpos30_7 in30 sp7 11140.846016
Rwpos30_8 in30 sp8 11140.846016
Rwpos30_9 in30 sp9 11140.846016
Rwpos30_10 in30 sp10 3183.098862
Rwpos30_11 in30 sp11 3183.098862
Rwpos30_12 in30 sp12 11140.846016
Rwpos30_13 in30 sp13 11140.846016
Rwpos30_14 in30 sp14 3183.098862
Rwpos30_15 in30 sp15 11140.846016
Rwpos30_16 in30 sp16 11140.846016
Rwpos30_17 in30 sp17 3183.098862
Rwpos30_18 in30 sp18 11140.846016
Rwpos30_19 in30 sp19 3183.098862
Rwpos30_20 in30 sp20 3183.098862
Rwpos30_21 in30 sp21 11140.846016
Rwpos30_22 in30 sp22 3183.098862
Rwpos30_23 in30 sp23 11140.846016
Rwpos30_24 in30 sp24 3183.098862
Rwpos30_25 in30 sp25 3183.098862
Rwpos30_26 in30 sp26 11140.846016
Rwpos30_27 in30 sp27 3183.098862
Rwpos30_28 in30 sp28 3183.098862
Rwpos30_29 in30 sp29 11140.846016
Rwpos30_30 in30 sp30 3183.098862
Rwpos30_31 in30 sp31 11140.846016
Rwpos30_32 in30 sp32 3183.098862
Rwpos30_33 in30 sp33 3183.098862
Rwpos30_34 in30 sp34 3183.098862
Rwpos30_35 in30 sp35 3183.098862
Rwpos30_36 in30 sp36 11140.846016
Rwpos30_37 in30 sp37 11140.846016
Rwpos30_38 in30 sp38 3183.098862
Rwpos30_39 in30 sp39 11140.846016
Rwpos30_40 in30 sp40 11140.846016
Rwpos30_41 in30 sp41 11140.846016
Rwpos30_42 in30 sp42 3183.098862
Rwpos30_43 in30 sp43 11140.846016
Rwpos30_44 in30 sp44 11140.846016
Rwpos30_45 in30 sp45 11140.846016
Rwpos30_46 in30 sp46 3183.098862
Rwpos30_47 in30 sp47 11140.846016
Rwpos30_48 in30 sp48 3183.098862
Rwpos30_49 in30 sp49 3183.098862
Rwpos30_50 in30 sp50 11140.846016
Rwpos30_51 in30 sp51 3183.098862
Rwpos30_52 in30 sp52 3183.098862
Rwpos30_53 in30 sp53 3183.098862
Rwpos30_54 in30 sp54 3183.098862
Rwpos30_55 in30 sp55 11140.846016
Rwpos30_56 in30 sp56 11140.846016
Rwpos30_57 in30 sp57 3183.098862
Rwpos30_58 in30 sp58 11140.846016
Rwpos30_59 in30 sp59 11140.846016
Rwpos30_60 in30 sp60 3183.098862
Rwpos30_61 in30 sp61 3183.098862
Rwpos30_62 in30 sp62 3183.098862
Rwpos30_63 in30 sp63 11140.846016
Rwpos30_64 in30 sp64 3183.098862
Rwpos30_65 in30 sp65 11140.846016
Rwpos30_66 in30 sp66 11140.846016
Rwpos30_67 in30 sp67 3183.098862
Rwpos30_68 in30 sp68 11140.846016
Rwpos30_69 in30 sp69 3183.098862
Rwpos30_70 in30 sp70 3183.098862
Rwpos30_71 in30 sp71 11140.846016
Rwpos30_72 in30 sp72 11140.846016
Rwpos30_73 in30 sp73 11140.846016
Rwpos30_74 in30 sp74 11140.846016
Rwpos30_75 in30 sp75 11140.846016
Rwpos30_76 in30 sp76 3183.098862
Rwpos30_77 in30 sp77 11140.846016
Rwpos30_78 in30 sp78 3183.098862
Rwpos30_79 in30 sp79 11140.846016
Rwpos30_80 in30 sp80 3183.098862
Rwpos30_81 in30 sp81 11140.846016
Rwpos30_82 in30 sp82 11140.846016
Rwpos30_83 in30 sp83 3183.098862
Rwpos30_84 in30 sp84 3183.098862
Rwpos30_85 in30 sp85 3183.098862
Rwpos30_86 in30 sp86 3183.098862
Rwpos30_87 in30 sp87 11140.846016
Rwpos30_88 in30 sp88 3183.098862
Rwpos30_89 in30 sp89 3183.098862
Rwpos30_90 in30 sp90 3183.098862
Rwpos30_91 in30 sp91 3183.098862
Rwpos30_92 in30 sp92 3183.098862
Rwpos30_93 in30 sp93 3183.098862
Rwpos30_94 in30 sp94 11140.846016
Rwpos30_95 in30 sp95 11140.846016
Rwpos30_96 in30 sp96 11140.846016
Rwpos30_97 in30 sp97 3183.098862
Rwpos30_98 in30 sp98 3183.098862
Rwpos30_99 in30 sp99 11140.846016
Rwpos30_100 in30 sp100 3183.098862
Rwpos31_1 in31 sp1 3183.098862
Rwpos31_2 in31 sp2 11140.846016
Rwpos31_3 in31 sp3 11140.846016
Rwpos31_4 in31 sp4 11140.846016
Rwpos31_5 in31 sp5 11140.846016
Rwpos31_6 in31 sp6 11140.846016
Rwpos31_7 in31 sp7 11140.846016
Rwpos31_8 in31 sp8 3183.098862
Rwpos31_9 in31 sp9 3183.098862
Rwpos31_10 in31 sp10 11140.846016
Rwpos31_11 in31 sp11 3183.098862
Rwpos31_12 in31 sp12 3183.098862
Rwpos31_13 in31 sp13 11140.846016
Rwpos31_14 in31 sp14 3183.098862
Rwpos31_15 in31 sp15 11140.846016
Rwpos31_16 in31 sp16 3183.098862
Rwpos31_17 in31 sp17 3183.098862
Rwpos31_18 in31 sp18 11140.846016
Rwpos31_19 in31 sp19 3183.098862
Rwpos31_20 in31 sp20 3183.098862
Rwpos31_21 in31 sp21 3183.098862
Rwpos31_22 in31 sp22 11140.846016
Rwpos31_23 in31 sp23 3183.098862
Rwpos31_24 in31 sp24 3183.098862
Rwpos31_25 in31 sp25 11140.846016
Rwpos31_26 in31 sp26 11140.846016
Rwpos31_27 in31 sp27 3183.098862
Rwpos31_28 in31 sp28 3183.098862
Rwpos31_29 in31 sp29 11140.846016
Rwpos31_30 in31 sp30 3183.098862
Rwpos31_31 in31 sp31 11140.846016
Rwpos31_32 in31 sp32 11140.846016
Rwpos31_33 in31 sp33 11140.846016
Rwpos31_34 in31 sp34 3183.098862
Rwpos31_35 in31 sp35 3183.098862
Rwpos31_36 in31 sp36 11140.846016
Rwpos31_37 in31 sp37 3183.098862
Rwpos31_38 in31 sp38 3183.098862
Rwpos31_39 in31 sp39 11140.846016
Rwpos31_40 in31 sp40 3183.098862
Rwpos31_41 in31 sp41 3183.098862
Rwpos31_42 in31 sp42 11140.846016
Rwpos31_43 in31 sp43 3183.098862
Rwpos31_44 in31 sp44 11140.846016
Rwpos31_45 in31 sp45 3183.098862
Rwpos31_46 in31 sp46 3183.098862
Rwpos31_47 in31 sp47 11140.846016
Rwpos31_48 in31 sp48 3183.098862
Rwpos31_49 in31 sp49 11140.846016
Rwpos31_50 in31 sp50 11140.846016
Rwpos31_51 in31 sp51 3183.098862
Rwpos31_52 in31 sp52 11140.846016
Rwpos31_53 in31 sp53 11140.846016
Rwpos31_54 in31 sp54 3183.098862
Rwpos31_55 in31 sp55 3183.098862
Rwpos31_56 in31 sp56 3183.098862
Rwpos31_57 in31 sp57 3183.098862
Rwpos31_58 in31 sp58 11140.846016
Rwpos31_59 in31 sp59 3183.098862
Rwpos31_60 in31 sp60 3183.098862
Rwpos31_61 in31 sp61 3183.098862
Rwpos31_62 in31 sp62 3183.098862
Rwpos31_63 in31 sp63 11140.846016
Rwpos31_64 in31 sp64 11140.846016
Rwpos31_65 in31 sp65 11140.846016
Rwpos31_66 in31 sp66 11140.846016
Rwpos31_67 in31 sp67 3183.098862
Rwpos31_68 in31 sp68 3183.098862
Rwpos31_69 in31 sp69 11140.846016
Rwpos31_70 in31 sp70 3183.098862
Rwpos31_71 in31 sp71 11140.846016
Rwpos31_72 in31 sp72 3183.098862
Rwpos31_73 in31 sp73 3183.098862
Rwpos31_74 in31 sp74 3183.098862
Rwpos31_75 in31 sp75 3183.098862
Rwpos31_76 in31 sp76 3183.098862
Rwpos31_77 in31 sp77 3183.098862
Rwpos31_78 in31 sp78 3183.098862
Rwpos31_79 in31 sp79 11140.846016
Rwpos31_80 in31 sp80 3183.098862
Rwpos31_81 in31 sp81 11140.846016
Rwpos31_82 in31 sp82 3183.098862
Rwpos31_83 in31 sp83 11140.846016
Rwpos31_84 in31 sp84 3183.098862
Rwpos31_85 in31 sp85 11140.846016
Rwpos31_86 in31 sp86 3183.098862
Rwpos31_87 in31 sp87 3183.098862
Rwpos31_88 in31 sp88 3183.098862
Rwpos31_89 in31 sp89 11140.846016
Rwpos31_90 in31 sp90 3183.098862
Rwpos31_91 in31 sp91 3183.098862
Rwpos31_92 in31 sp92 3183.098862
Rwpos31_93 in31 sp93 11140.846016
Rwpos31_94 in31 sp94 11140.846016
Rwpos31_95 in31 sp95 11140.846016
Rwpos31_96 in31 sp96 11140.846016
Rwpos31_97 in31 sp97 3183.098862
Rwpos31_98 in31 sp98 3183.098862
Rwpos31_99 in31 sp99 11140.846016
Rwpos31_100 in31 sp100 3183.098862
Rwpos32_1 in32 sp1 11140.846016
Rwpos32_2 in32 sp2 3183.098862
Rwpos32_3 in32 sp3 3183.098862
Rwpos32_4 in32 sp4 11140.846016
Rwpos32_5 in32 sp5 11140.846016
Rwpos32_6 in32 sp6 11140.846016
Rwpos32_7 in32 sp7 3183.098862
Rwpos32_8 in32 sp8 3183.098862
Rwpos32_9 in32 sp9 3183.098862
Rwpos32_10 in32 sp10 3183.098862
Rwpos32_11 in32 sp11 11140.846016
Rwpos32_12 in32 sp12 11140.846016
Rwpos32_13 in32 sp13 3183.098862
Rwpos32_14 in32 sp14 3183.098862
Rwpos32_15 in32 sp15 11140.846016
Rwpos32_16 in32 sp16 3183.098862
Rwpos32_17 in32 sp17 11140.846016
Rwpos32_18 in32 sp18 3183.098862
Rwpos32_19 in32 sp19 3183.098862
Rwpos32_20 in32 sp20 11140.846016
Rwpos32_21 in32 sp21 3183.098862
Rwpos32_22 in32 sp22 3183.098862
Rwpos32_23 in32 sp23 3183.098862
Rwpos32_24 in32 sp24 11140.846016
Rwpos32_25 in32 sp25 11140.846016
Rwpos32_26 in32 sp26 11140.846016
Rwpos32_27 in32 sp27 11140.846016
Rwpos32_28 in32 sp28 3183.098862
Rwpos32_29 in32 sp29 3183.098862
Rwpos32_30 in32 sp30 3183.098862
Rwpos32_31 in32 sp31 3183.098862
Rwpos32_32 in32 sp32 11140.846016
Rwpos32_33 in32 sp33 3183.098862
Rwpos32_34 in32 sp34 11140.846016
Rwpos32_35 in32 sp35 11140.846016
Rwpos32_36 in32 sp36 3183.098862
Rwpos32_37 in32 sp37 3183.098862
Rwpos32_38 in32 sp38 11140.846016
Rwpos32_39 in32 sp39 3183.098862
Rwpos32_40 in32 sp40 3183.098862
Rwpos32_41 in32 sp41 3183.098862
Rwpos32_42 in32 sp42 3183.098862
Rwpos32_43 in32 sp43 3183.098862
Rwpos32_44 in32 sp44 3183.098862
Rwpos32_45 in32 sp45 11140.846016
Rwpos32_46 in32 sp46 11140.846016
Rwpos32_47 in32 sp47 3183.098862
Rwpos32_48 in32 sp48 3183.098862
Rwpos32_49 in32 sp49 11140.846016
Rwpos32_50 in32 sp50 11140.846016
Rwpos32_51 in32 sp51 11140.846016
Rwpos32_52 in32 sp52 11140.846016
Rwpos32_53 in32 sp53 3183.098862
Rwpos32_54 in32 sp54 3183.098862
Rwpos32_55 in32 sp55 3183.098862
Rwpos32_56 in32 sp56 3183.098862
Rwpos32_57 in32 sp57 11140.846016
Rwpos32_58 in32 sp58 11140.846016
Rwpos32_59 in32 sp59 3183.098862
Rwpos32_60 in32 sp60 11140.846016
Rwpos32_61 in32 sp61 11140.846016
Rwpos32_62 in32 sp62 3183.098862
Rwpos32_63 in32 sp63 11140.846016
Rwpos32_64 in32 sp64 3183.098862
Rwpos32_65 in32 sp65 11140.846016
Rwpos32_66 in32 sp66 3183.098862
Rwpos32_67 in32 sp67 3183.098862
Rwpos32_68 in32 sp68 3183.098862
Rwpos32_69 in32 sp69 3183.098862
Rwpos32_70 in32 sp70 11140.846016
Rwpos32_71 in32 sp71 11140.846016
Rwpos32_72 in32 sp72 11140.846016
Rwpos32_73 in32 sp73 11140.846016
Rwpos32_74 in32 sp74 3183.098862
Rwpos32_75 in32 sp75 3183.098862
Rwpos32_76 in32 sp76 11140.846016
Rwpos32_77 in32 sp77 3183.098862
Rwpos32_78 in32 sp78 11140.846016
Rwpos32_79 in32 sp79 11140.846016
Rwpos32_80 in32 sp80 3183.098862
Rwpos32_81 in32 sp81 11140.846016
Rwpos32_82 in32 sp82 3183.098862
Rwpos32_83 in32 sp83 3183.098862
Rwpos32_84 in32 sp84 3183.098862
Rwpos32_85 in32 sp85 11140.846016
Rwpos32_86 in32 sp86 11140.846016
Rwpos32_87 in32 sp87 3183.098862
Rwpos32_88 in32 sp88 3183.098862
Rwpos32_89 in32 sp89 11140.846016
Rwpos32_90 in32 sp90 11140.846016
Rwpos32_91 in32 sp91 3183.098862
Rwpos32_92 in32 sp92 11140.846016
Rwpos32_93 in32 sp93 3183.098862
Rwpos32_94 in32 sp94 3183.098862
Rwpos32_95 in32 sp95 11140.846016
Rwpos32_96 in32 sp96 11140.846016
Rwpos32_97 in32 sp97 11140.846016
Rwpos32_98 in32 sp98 3183.098862
Rwpos32_99 in32 sp99 3183.098862
Rwpos32_100 in32 sp100 11140.846016
Rwpos33_1 in33 sp1 11140.846016
Rwpos33_2 in33 sp2 3183.098862
Rwpos33_3 in33 sp3 11140.846016
Rwpos33_4 in33 sp4 11140.846016
Rwpos33_5 in33 sp5 3183.098862
Rwpos33_6 in33 sp6 11140.846016
Rwpos33_7 in33 sp7 3183.098862
Rwpos33_8 in33 sp8 3183.098862
Rwpos33_9 in33 sp9 3183.098862
Rwpos33_10 in33 sp10 3183.098862
Rwpos33_11 in33 sp11 11140.846016
Rwpos33_12 in33 sp12 3183.098862
Rwpos33_13 in33 sp13 11140.846016
Rwpos33_14 in33 sp14 3183.098862
Rwpos33_15 in33 sp15 11140.846016
Rwpos33_16 in33 sp16 3183.098862
Rwpos33_17 in33 sp17 11140.846016
Rwpos33_18 in33 sp18 11140.846016
Rwpos33_19 in33 sp19 3183.098862
Rwpos33_20 in33 sp20 11140.846016
Rwpos33_21 in33 sp21 11140.846016
Rwpos33_22 in33 sp22 3183.098862
Rwpos33_23 in33 sp23 3183.098862
Rwpos33_24 in33 sp24 3183.098862
Rwpos33_25 in33 sp25 3183.098862
Rwpos33_26 in33 sp26 11140.846016
Rwpos33_27 in33 sp27 11140.846016
Rwpos33_28 in33 sp28 3183.098862
Rwpos33_29 in33 sp29 11140.846016
Rwpos33_30 in33 sp30 3183.098862
Rwpos33_31 in33 sp31 11140.846016
Rwpos33_32 in33 sp32 3183.098862
Rwpos33_33 in33 sp33 11140.846016
Rwpos33_34 in33 sp34 11140.846016
Rwpos33_35 in33 sp35 3183.098862
Rwpos33_36 in33 sp36 11140.846016
Rwpos33_37 in33 sp37 11140.846016
Rwpos33_38 in33 sp38 11140.846016
Rwpos33_39 in33 sp39 11140.846016
Rwpos33_40 in33 sp40 3183.098862
Rwpos33_41 in33 sp41 11140.846016
Rwpos33_42 in33 sp42 11140.846016
Rwpos33_43 in33 sp43 11140.846016
Rwpos33_44 in33 sp44 11140.846016
Rwpos33_45 in33 sp45 11140.846016
Rwpos33_46 in33 sp46 11140.846016
Rwpos33_47 in33 sp47 11140.846016
Rwpos33_48 in33 sp48 3183.098862
Rwpos33_49 in33 sp49 11140.846016
Rwpos33_50 in33 sp50 3183.098862
Rwpos33_51 in33 sp51 3183.098862
Rwpos33_52 in33 sp52 11140.846016
Rwpos33_53 in33 sp53 11140.846016
Rwpos33_54 in33 sp54 11140.846016
Rwpos33_55 in33 sp55 3183.098862
Rwpos33_56 in33 sp56 11140.846016
Rwpos33_57 in33 sp57 3183.098862
Rwpos33_58 in33 sp58 11140.846016
Rwpos33_59 in33 sp59 11140.846016
Rwpos33_60 in33 sp60 3183.098862
Rwpos33_61 in33 sp61 3183.098862
Rwpos33_62 in33 sp62 3183.098862
Rwpos33_63 in33 sp63 11140.846016
Rwpos33_64 in33 sp64 3183.098862
Rwpos33_65 in33 sp65 11140.846016
Rwpos33_66 in33 sp66 11140.846016
Rwpos33_67 in33 sp67 3183.098862
Rwpos33_68 in33 sp68 11140.846016
Rwpos33_69 in33 sp69 3183.098862
Rwpos33_70 in33 sp70 3183.098862
Rwpos33_71 in33 sp71 3183.098862
Rwpos33_72 in33 sp72 3183.098862
Rwpos33_73 in33 sp73 3183.098862
Rwpos33_74 in33 sp74 3183.098862
Rwpos33_75 in33 sp75 11140.846016
Rwpos33_76 in33 sp76 11140.846016
Rwpos33_77 in33 sp77 3183.098862
Rwpos33_78 in33 sp78 3183.098862
Rwpos33_79 in33 sp79 3183.098862
Rwpos33_80 in33 sp80 11140.846016
Rwpos33_81 in33 sp81 11140.846016
Rwpos33_82 in33 sp82 11140.846016
Rwpos33_83 in33 sp83 3183.098862
Rwpos33_84 in33 sp84 3183.098862
Rwpos33_85 in33 sp85 11140.846016
Rwpos33_86 in33 sp86 11140.846016
Rwpos33_87 in33 sp87 3183.098862
Rwpos33_88 in33 sp88 11140.846016
Rwpos33_89 in33 sp89 11140.846016
Rwpos33_90 in33 sp90 3183.098862
Rwpos33_91 in33 sp91 11140.846016
Rwpos33_92 in33 sp92 3183.098862
Rwpos33_93 in33 sp93 3183.098862
Rwpos33_94 in33 sp94 3183.098862
Rwpos33_95 in33 sp95 11140.846016
Rwpos33_96 in33 sp96 3183.098862
Rwpos33_97 in33 sp97 11140.846016
Rwpos33_98 in33 sp98 11140.846016
Rwpos33_99 in33 sp99 3183.098862
Rwpos33_100 in33 sp100 11140.846016
Rwpos34_1 in34 sp1 3183.098862
Rwpos34_2 in34 sp2 3183.098862
Rwpos34_3 in34 sp3 3183.098862
Rwpos34_4 in34 sp4 3183.098862
Rwpos34_5 in34 sp5 11140.846016
Rwpos34_6 in34 sp6 11140.846016
Rwpos34_7 in34 sp7 11140.846016
Rwpos34_8 in34 sp8 11140.846016
Rwpos34_9 in34 sp9 11140.846016
Rwpos34_10 in34 sp10 11140.846016
Rwpos34_11 in34 sp11 11140.846016
Rwpos34_12 in34 sp12 11140.846016
Rwpos34_13 in34 sp13 3183.098862
Rwpos34_14 in34 sp14 3183.098862
Rwpos34_15 in34 sp15 11140.846016
Rwpos34_16 in34 sp16 11140.846016
Rwpos34_17 in34 sp17 3183.098862
Rwpos34_18 in34 sp18 3183.098862
Rwpos34_19 in34 sp19 3183.098862
Rwpos34_20 in34 sp20 3183.098862
Rwpos34_21 in34 sp21 11140.846016
Rwpos34_22 in34 sp22 3183.098862
Rwpos34_23 in34 sp23 11140.846016
Rwpos34_24 in34 sp24 3183.098862
Rwpos34_25 in34 sp25 11140.846016
Rwpos34_26 in34 sp26 3183.098862
Rwpos34_27 in34 sp27 11140.846016
Rwpos34_28 in34 sp28 11140.846016
Rwpos34_29 in34 sp29 11140.846016
Rwpos34_30 in34 sp30 3183.098862
Rwpos34_31 in34 sp31 11140.846016
Rwpos34_32 in34 sp32 3183.098862
Rwpos34_33 in34 sp33 3183.098862
Rwpos34_34 in34 sp34 3183.098862
Rwpos34_35 in34 sp35 11140.846016
Rwpos34_36 in34 sp36 11140.846016
Rwpos34_37 in34 sp37 11140.846016
Rwpos34_38 in34 sp38 3183.098862
Rwpos34_39 in34 sp39 3183.098862
Rwpos34_40 in34 sp40 11140.846016
Rwpos34_41 in34 sp41 3183.098862
Rwpos34_42 in34 sp42 11140.846016
Rwpos34_43 in34 sp43 11140.846016
Rwpos34_44 in34 sp44 3183.098862
Rwpos34_45 in34 sp45 11140.846016
Rwpos34_46 in34 sp46 3183.098862
Rwpos34_47 in34 sp47 11140.846016
Rwpos34_48 in34 sp48 3183.098862
Rwpos34_49 in34 sp49 3183.098862
Rwpos34_50 in34 sp50 3183.098862
Rwpos34_51 in34 sp51 3183.098862
Rwpos34_52 in34 sp52 11140.846016
Rwpos34_53 in34 sp53 3183.098862
Rwpos34_54 in34 sp54 3183.098862
Rwpos34_55 in34 sp55 11140.846016
Rwpos34_56 in34 sp56 11140.846016
Rwpos34_57 in34 sp57 3183.098862
Rwpos34_58 in34 sp58 11140.846016
Rwpos34_59 in34 sp59 11140.846016
Rwpos34_60 in34 sp60 3183.098862
Rwpos34_61 in34 sp61 3183.098862
Rwpos34_62 in34 sp62 3183.098862
Rwpos34_63 in34 sp63 11140.846016
Rwpos34_64 in34 sp64 3183.098862
Rwpos34_65 in34 sp65 3183.098862
Rwpos34_66 in34 sp66 11140.846016
Rwpos34_67 in34 sp67 11140.846016
Rwpos34_68 in34 sp68 11140.846016
Rwpos34_69 in34 sp69 3183.098862
Rwpos34_70 in34 sp70 3183.098862
Rwpos34_71 in34 sp71 11140.846016
Rwpos34_72 in34 sp72 11140.846016
Rwpos34_73 in34 sp73 11140.846016
Rwpos34_74 in34 sp74 3183.098862
Rwpos34_75 in34 sp75 3183.098862
Rwpos34_76 in34 sp76 11140.846016
Rwpos34_77 in34 sp77 3183.098862
Rwpos34_78 in34 sp78 3183.098862
Rwpos34_79 in34 sp79 11140.846016
Rwpos34_80 in34 sp80 3183.098862
Rwpos34_81 in34 sp81 3183.098862
Rwpos34_82 in34 sp82 3183.098862
Rwpos34_83 in34 sp83 3183.098862
Rwpos34_84 in34 sp84 3183.098862
Rwpos34_85 in34 sp85 11140.846016
Rwpos34_86 in34 sp86 3183.098862
Rwpos34_87 in34 sp87 11140.846016
Rwpos34_88 in34 sp88 11140.846016
Rwpos34_89 in34 sp89 3183.098862
Rwpos34_90 in34 sp90 11140.846016
Rwpos34_91 in34 sp91 3183.098862
Rwpos34_92 in34 sp92 3183.098862
Rwpos34_93 in34 sp93 3183.098862
Rwpos34_94 in34 sp94 3183.098862
Rwpos34_95 in34 sp95 11140.846016
Rwpos34_96 in34 sp96 3183.098862
Rwpos34_97 in34 sp97 3183.098862
Rwpos34_98 in34 sp98 11140.846016
Rwpos34_99 in34 sp99 3183.098862
Rwpos34_100 in34 sp100 11140.846016
Rwpos35_1 in35 sp1 11140.846016
Rwpos35_2 in35 sp2 3183.098862
Rwpos35_3 in35 sp3 3183.098862
Rwpos35_4 in35 sp4 3183.098862
Rwpos35_5 in35 sp5 11140.846016
Rwpos35_6 in35 sp6 11140.846016
Rwpos35_7 in35 sp7 3183.098862
Rwpos35_8 in35 sp8 11140.846016
Rwpos35_9 in35 sp9 11140.846016
Rwpos35_10 in35 sp10 3183.098862
Rwpos35_11 in35 sp11 11140.846016
Rwpos35_12 in35 sp12 11140.846016
Rwpos35_13 in35 sp13 11140.846016
Rwpos35_14 in35 sp14 3183.098862
Rwpos35_15 in35 sp15 11140.846016
Rwpos35_16 in35 sp16 3183.098862
Rwpos35_17 in35 sp17 11140.846016
Rwpos35_18 in35 sp18 3183.098862
Rwpos35_19 in35 sp19 11140.846016
Rwpos35_20 in35 sp20 11140.846016
Rwpos35_21 in35 sp21 3183.098862
Rwpos35_22 in35 sp22 3183.098862
Rwpos35_23 in35 sp23 11140.846016
Rwpos35_24 in35 sp24 3183.098862
Rwpos35_25 in35 sp25 3183.098862
Rwpos35_26 in35 sp26 3183.098862
Rwpos35_27 in35 sp27 11140.846016
Rwpos35_28 in35 sp28 3183.098862
Rwpos35_29 in35 sp29 3183.098862
Rwpos35_30 in35 sp30 3183.098862
Rwpos35_31 in35 sp31 3183.098862
Rwpos35_32 in35 sp32 3183.098862
Rwpos35_33 in35 sp33 11140.846016
Rwpos35_34 in35 sp34 3183.098862
Rwpos35_35 in35 sp35 3183.098862
Rwpos35_36 in35 sp36 11140.846016
Rwpos35_37 in35 sp37 11140.846016
Rwpos35_38 in35 sp38 11140.846016
Rwpos35_39 in35 sp39 11140.846016
Rwpos35_40 in35 sp40 3183.098862
Rwpos35_41 in35 sp41 3183.098862
Rwpos35_42 in35 sp42 3183.098862
Rwpos35_43 in35 sp43 3183.098862
Rwpos35_44 in35 sp44 11140.846016
Rwpos35_45 in35 sp45 11140.846016
Rwpos35_46 in35 sp46 3183.098862
Rwpos35_47 in35 sp47 11140.846016
Rwpos35_48 in35 sp48 11140.846016
Rwpos35_49 in35 sp49 11140.846016
Rwpos35_50 in35 sp50 3183.098862
Rwpos35_51 in35 sp51 3183.098862
Rwpos35_52 in35 sp52 11140.846016
Rwpos35_53 in35 sp53 3183.098862
Rwpos35_54 in35 sp54 3183.098862
Rwpos35_55 in35 sp55 3183.098862
Rwpos35_56 in35 sp56 3183.098862
Rwpos35_57 in35 sp57 11140.846016
Rwpos35_58 in35 sp58 11140.846016
Rwpos35_59 in35 sp59 11140.846016
Rwpos35_60 in35 sp60 11140.846016
Rwpos35_61 in35 sp61 11140.846016
Rwpos35_62 in35 sp62 3183.098862
Rwpos35_63 in35 sp63 11140.846016
Rwpos35_64 in35 sp64 11140.846016
Rwpos35_65 in35 sp65 3183.098862
Rwpos35_66 in35 sp66 3183.098862
Rwpos35_67 in35 sp67 11140.846016
Rwpos35_68 in35 sp68 11140.846016
Rwpos35_69 in35 sp69 11140.846016
Rwpos35_70 in35 sp70 11140.846016
Rwpos35_71 in35 sp71 11140.846016
Rwpos35_72 in35 sp72 3183.098862
Rwpos35_73 in35 sp73 3183.098862
Rwpos35_74 in35 sp74 11140.846016
Rwpos35_75 in35 sp75 3183.098862
Rwpos35_76 in35 sp76 11140.846016
Rwpos35_77 in35 sp77 3183.098862
Rwpos35_78 in35 sp78 3183.098862
Rwpos35_79 in35 sp79 11140.846016
Rwpos35_80 in35 sp80 3183.098862
Rwpos35_81 in35 sp81 11140.846016
Rwpos35_82 in35 sp82 11140.846016
Rwpos35_83 in35 sp83 3183.098862
Rwpos35_84 in35 sp84 11140.846016
Rwpos35_85 in35 sp85 11140.846016
Rwpos35_86 in35 sp86 11140.846016
Rwpos35_87 in35 sp87 3183.098862
Rwpos35_88 in35 sp88 3183.098862
Rwpos35_89 in35 sp89 3183.098862
Rwpos35_90 in35 sp90 11140.846016
Rwpos35_91 in35 sp91 3183.098862
Rwpos35_92 in35 sp92 3183.098862
Rwpos35_93 in35 sp93 3183.098862
Rwpos35_94 in35 sp94 3183.098862
Rwpos35_95 in35 sp95 3183.098862
Rwpos35_96 in35 sp96 11140.846016
Rwpos35_97 in35 sp97 3183.098862
Rwpos35_98 in35 sp98 11140.846016
Rwpos35_99 in35 sp99 11140.846016
Rwpos35_100 in35 sp100 3183.098862
Rwpos36_1 in36 sp1 11140.846016
Rwpos36_2 in36 sp2 11140.846016
Rwpos36_3 in36 sp3 11140.846016
Rwpos36_4 in36 sp4 3183.098862
Rwpos36_5 in36 sp5 3183.098862
Rwpos36_6 in36 sp6 11140.846016
Rwpos36_7 in36 sp7 3183.098862
Rwpos36_8 in36 sp8 3183.098862
Rwpos36_9 in36 sp9 3183.098862
Rwpos36_10 in36 sp10 3183.098862
Rwpos36_11 in36 sp11 11140.846016
Rwpos36_12 in36 sp12 3183.098862
Rwpos36_13 in36 sp13 11140.846016
Rwpos36_14 in36 sp14 11140.846016
Rwpos36_15 in36 sp15 3183.098862
Rwpos36_16 in36 sp16 3183.098862
Rwpos36_17 in36 sp17 11140.846016
Rwpos36_18 in36 sp18 11140.846016
Rwpos36_19 in36 sp19 3183.098862
Rwpos36_20 in36 sp20 3183.098862
Rwpos36_21 in36 sp21 3183.098862
Rwpos36_22 in36 sp22 3183.098862
Rwpos36_23 in36 sp23 3183.098862
Rwpos36_24 in36 sp24 3183.098862
Rwpos36_25 in36 sp25 3183.098862
Rwpos36_26 in36 sp26 3183.098862
Rwpos36_27 in36 sp27 11140.846016
Rwpos36_28 in36 sp28 3183.098862
Rwpos36_29 in36 sp29 11140.846016
Rwpos36_30 in36 sp30 11140.846016
Rwpos36_31 in36 sp31 3183.098862
Rwpos36_32 in36 sp32 3183.098862
Rwpos36_33 in36 sp33 11140.846016
Rwpos36_34 in36 sp34 3183.098862
Rwpos36_35 in36 sp35 3183.098862
Rwpos36_36 in36 sp36 3183.098862
Rwpos36_37 in36 sp37 3183.098862
Rwpos36_38 in36 sp38 11140.846016
Rwpos36_39 in36 sp39 11140.846016
Rwpos36_40 in36 sp40 3183.098862
Rwpos36_41 in36 sp41 11140.846016
Rwpos36_42 in36 sp42 11140.846016
Rwpos36_43 in36 sp43 11140.846016
Rwpos36_44 in36 sp44 3183.098862
Rwpos36_45 in36 sp45 3183.098862
Rwpos36_46 in36 sp46 3183.098862
Rwpos36_47 in36 sp47 11140.846016
Rwpos36_48 in36 sp48 11140.846016
Rwpos36_49 in36 sp49 11140.846016
Rwpos36_50 in36 sp50 11140.846016
Rwpos36_51 in36 sp51 3183.098862
Rwpos36_52 in36 sp52 11140.846016
Rwpos36_53 in36 sp53 3183.098862
Rwpos36_54 in36 sp54 3183.098862
Rwpos36_55 in36 sp55 11140.846016
Rwpos36_56 in36 sp56 3183.098862
Rwpos36_57 in36 sp57 3183.098862
Rwpos36_58 in36 sp58 3183.098862
Rwpos36_59 in36 sp59 3183.098862
Rwpos36_60 in36 sp60 3183.098862
Rwpos36_61 in36 sp61 11140.846016
Rwpos36_62 in36 sp62 3183.098862
Rwpos36_63 in36 sp63 3183.098862
Rwpos36_64 in36 sp64 3183.098862
Rwpos36_65 in36 sp65 11140.846016
Rwpos36_66 in36 sp66 3183.098862
Rwpos36_67 in36 sp67 11140.846016
Rwpos36_68 in36 sp68 3183.098862
Rwpos36_69 in36 sp69 11140.846016
Rwpos36_70 in36 sp70 11140.846016
Rwpos36_71 in36 sp71 3183.098862
Rwpos36_72 in36 sp72 3183.098862
Rwpos36_73 in36 sp73 3183.098862
Rwpos36_74 in36 sp74 11140.846016
Rwpos36_75 in36 sp75 3183.098862
Rwpos36_76 in36 sp76 11140.846016
Rwpos36_77 in36 sp77 3183.098862
Rwpos36_78 in36 sp78 3183.098862
Rwpos36_79 in36 sp79 3183.098862
Rwpos36_80 in36 sp80 3183.098862
Rwpos36_81 in36 sp81 11140.846016
Rwpos36_82 in36 sp82 3183.098862
Rwpos36_83 in36 sp83 3183.098862
Rwpos36_84 in36 sp84 3183.098862
Rwpos36_85 in36 sp85 3183.098862
Rwpos36_86 in36 sp86 3183.098862
Rwpos36_87 in36 sp87 11140.846016
Rwpos36_88 in36 sp88 11140.846016
Rwpos36_89 in36 sp89 11140.846016
Rwpos36_90 in36 sp90 11140.846016
Rwpos36_91 in36 sp91 3183.098862
Rwpos36_92 in36 sp92 3183.098862
Rwpos36_93 in36 sp93 3183.098862
Rwpos36_94 in36 sp94 3183.098862
Rwpos36_95 in36 sp95 11140.846016
Rwpos36_96 in36 sp96 3183.098862
Rwpos36_97 in36 sp97 3183.098862
Rwpos36_98 in36 sp98 11140.846016
Rwpos36_99 in36 sp99 11140.846016
Rwpos36_100 in36 sp100 11140.846016
Rwpos37_1 in37 sp1 3183.098862
Rwpos37_2 in37 sp2 3183.098862
Rwpos37_3 in37 sp3 11140.846016
Rwpos37_4 in37 sp4 11140.846016
Rwpos37_5 in37 sp5 3183.098862
Rwpos37_6 in37 sp6 11140.846016
Rwpos37_7 in37 sp7 3183.098862
Rwpos37_8 in37 sp8 3183.098862
Rwpos37_9 in37 sp9 3183.098862
Rwpos37_10 in37 sp10 11140.846016
Rwpos37_11 in37 sp11 3183.098862
Rwpos37_12 in37 sp12 11140.846016
Rwpos37_13 in37 sp13 11140.846016
Rwpos37_14 in37 sp14 3183.098862
Rwpos37_15 in37 sp15 3183.098862
Rwpos37_16 in37 sp16 11140.846016
Rwpos37_17 in37 sp17 3183.098862
Rwpos37_18 in37 sp18 11140.846016
Rwpos37_19 in37 sp19 11140.846016
Rwpos37_20 in37 sp20 3183.098862
Rwpos37_21 in37 sp21 11140.846016
Rwpos37_22 in37 sp22 3183.098862
Rwpos37_23 in37 sp23 11140.846016
Rwpos37_24 in37 sp24 11140.846016
Rwpos37_25 in37 sp25 11140.846016
Rwpos37_26 in37 sp26 3183.098862
Rwpos37_27 in37 sp27 11140.846016
Rwpos37_28 in37 sp28 11140.846016
Rwpos37_29 in37 sp29 3183.098862
Rwpos37_30 in37 sp30 11140.846016
Rwpos37_31 in37 sp31 11140.846016
Rwpos37_32 in37 sp32 11140.846016
Rwpos37_33 in37 sp33 11140.846016
Rwpos37_34 in37 sp34 3183.098862
Rwpos37_35 in37 sp35 11140.846016
Rwpos37_36 in37 sp36 3183.098862
Rwpos37_37 in37 sp37 11140.846016
Rwpos37_38 in37 sp38 11140.846016
Rwpos37_39 in37 sp39 11140.846016
Rwpos37_40 in37 sp40 3183.098862
Rwpos37_41 in37 sp41 3183.098862
Rwpos37_42 in37 sp42 11140.846016
Rwpos37_43 in37 sp43 11140.846016
Rwpos37_44 in37 sp44 11140.846016
Rwpos37_45 in37 sp45 11140.846016
Rwpos37_46 in37 sp46 3183.098862
Rwpos37_47 in37 sp47 3183.098862
Rwpos37_48 in37 sp48 3183.098862
Rwpos37_49 in37 sp49 3183.098862
Rwpos37_50 in37 sp50 11140.846016
Rwpos37_51 in37 sp51 3183.098862
Rwpos37_52 in37 sp52 3183.098862
Rwpos37_53 in37 sp53 3183.098862
Rwpos37_54 in37 sp54 11140.846016
Rwpos37_55 in37 sp55 11140.846016
Rwpos37_56 in37 sp56 11140.846016
Rwpos37_57 in37 sp57 3183.098862
Rwpos37_58 in37 sp58 3183.098862
Rwpos37_59 in37 sp59 3183.098862
Rwpos37_60 in37 sp60 3183.098862
Rwpos37_61 in37 sp61 11140.846016
Rwpos37_62 in37 sp62 3183.098862
Rwpos37_63 in37 sp63 11140.846016
Rwpos37_64 in37 sp64 3183.098862
Rwpos37_65 in37 sp65 11140.846016
Rwpos37_66 in37 sp66 11140.846016
Rwpos37_67 in37 sp67 3183.098862
Rwpos37_68 in37 sp68 3183.098862
Rwpos37_69 in37 sp69 3183.098862
Rwpos37_70 in37 sp70 3183.098862
Rwpos37_71 in37 sp71 3183.098862
Rwpos37_72 in37 sp72 11140.846016
Rwpos37_73 in37 sp73 3183.098862
Rwpos37_74 in37 sp74 3183.098862
Rwpos37_75 in37 sp75 11140.846016
Rwpos37_76 in37 sp76 3183.098862
Rwpos37_77 in37 sp77 3183.098862
Rwpos37_78 in37 sp78 11140.846016
Rwpos37_79 in37 sp79 11140.846016
Rwpos37_80 in37 sp80 11140.846016
Rwpos37_81 in37 sp81 11140.846016
Rwpos37_82 in37 sp82 3183.098862
Rwpos37_83 in37 sp83 3183.098862
Rwpos37_84 in37 sp84 11140.846016
Rwpos37_85 in37 sp85 11140.846016
Rwpos37_86 in37 sp86 3183.098862
Rwpos37_87 in37 sp87 3183.098862
Rwpos37_88 in37 sp88 3183.098862
Rwpos37_89 in37 sp89 11140.846016
Rwpos37_90 in37 sp90 3183.098862
Rwpos37_91 in37 sp91 11140.846016
Rwpos37_92 in37 sp92 3183.098862
Rwpos37_93 in37 sp93 3183.098862
Rwpos37_94 in37 sp94 3183.098862
Rwpos37_95 in37 sp95 3183.098862
Rwpos37_96 in37 sp96 3183.098862
Rwpos37_97 in37 sp97 11140.846016
Rwpos37_98 in37 sp98 11140.846016
Rwpos37_99 in37 sp99 3183.098862
Rwpos37_100 in37 sp100 11140.846016
Rwpos38_1 in38 sp1 11140.846016
Rwpos38_2 in38 sp2 3183.098862
Rwpos38_3 in38 sp3 3183.098862
Rwpos38_4 in38 sp4 3183.098862
Rwpos38_5 in38 sp5 3183.098862
Rwpos38_6 in38 sp6 11140.846016
Rwpos38_7 in38 sp7 11140.846016
Rwpos38_8 in38 sp8 11140.846016
Rwpos38_9 in38 sp9 11140.846016
Rwpos38_10 in38 sp10 3183.098862
Rwpos38_11 in38 sp11 3183.098862
Rwpos38_12 in38 sp12 3183.098862
Rwpos38_13 in38 sp13 3183.098862
Rwpos38_14 in38 sp14 3183.098862
Rwpos38_15 in38 sp15 3183.098862
Rwpos38_16 in38 sp16 11140.846016
Rwpos38_17 in38 sp17 11140.846016
Rwpos38_18 in38 sp18 3183.098862
Rwpos38_19 in38 sp19 3183.098862
Rwpos38_20 in38 sp20 11140.846016
Rwpos38_21 in38 sp21 3183.098862
Rwpos38_22 in38 sp22 11140.846016
Rwpos38_23 in38 sp23 3183.098862
Rwpos38_24 in38 sp24 11140.846016
Rwpos38_25 in38 sp25 11140.846016
Rwpos38_26 in38 sp26 11140.846016
Rwpos38_27 in38 sp27 11140.846016
Rwpos38_28 in38 sp28 11140.846016
Rwpos38_29 in38 sp29 3183.098862
Rwpos38_30 in38 sp30 11140.846016
Rwpos38_31 in38 sp31 3183.098862
Rwpos38_32 in38 sp32 11140.846016
Rwpos38_33 in38 sp33 11140.846016
Rwpos38_34 in38 sp34 3183.098862
Rwpos38_35 in38 sp35 3183.098862
Rwpos38_36 in38 sp36 3183.098862
Rwpos38_37 in38 sp37 3183.098862
Rwpos38_38 in38 sp38 3183.098862
Rwpos38_39 in38 sp39 3183.098862
Rwpos38_40 in38 sp40 3183.098862
Rwpos38_41 in38 sp41 11140.846016
Rwpos38_42 in38 sp42 3183.098862
Rwpos38_43 in38 sp43 11140.846016
Rwpos38_44 in38 sp44 11140.846016
Rwpos38_45 in38 sp45 11140.846016
Rwpos38_46 in38 sp46 3183.098862
Rwpos38_47 in38 sp47 3183.098862
Rwpos38_48 in38 sp48 3183.098862
Rwpos38_49 in38 sp49 11140.846016
Rwpos38_50 in38 sp50 3183.098862
Rwpos38_51 in38 sp51 3183.098862
Rwpos38_52 in38 sp52 11140.846016
Rwpos38_53 in38 sp53 3183.098862
Rwpos38_54 in38 sp54 3183.098862
Rwpos38_55 in38 sp55 3183.098862
Rwpos38_56 in38 sp56 3183.098862
Rwpos38_57 in38 sp57 11140.846016
Rwpos38_58 in38 sp58 3183.098862
Rwpos38_59 in38 sp59 11140.846016
Rwpos38_60 in38 sp60 3183.098862
Rwpos38_61 in38 sp61 11140.846016
Rwpos38_62 in38 sp62 3183.098862
Rwpos38_63 in38 sp63 11140.846016
Rwpos38_64 in38 sp64 3183.098862
Rwpos38_65 in38 sp65 11140.846016
Rwpos38_66 in38 sp66 3183.098862
Rwpos38_67 in38 sp67 3183.098862
Rwpos38_68 in38 sp68 3183.098862
Rwpos38_69 in38 sp69 11140.846016
Rwpos38_70 in38 sp70 3183.098862
Rwpos38_71 in38 sp71 3183.098862
Rwpos38_72 in38 sp72 3183.098862
Rwpos38_73 in38 sp73 11140.846016
Rwpos38_74 in38 sp74 3183.098862
Rwpos38_75 in38 sp75 11140.846016
Rwpos38_76 in38 sp76 3183.098862
Rwpos38_77 in38 sp77 11140.846016
Rwpos38_78 in38 sp78 3183.098862
Rwpos38_79 in38 sp79 11140.846016
Rwpos38_80 in38 sp80 11140.846016
Rwpos38_81 in38 sp81 3183.098862
Rwpos38_82 in38 sp82 11140.846016
Rwpos38_83 in38 sp83 11140.846016
Rwpos38_84 in38 sp84 3183.098862
Rwpos38_85 in38 sp85 3183.098862
Rwpos38_86 in38 sp86 3183.098862
Rwpos38_87 in38 sp87 3183.098862
Rwpos38_88 in38 sp88 3183.098862
Rwpos38_89 in38 sp89 11140.846016
Rwpos38_90 in38 sp90 11140.846016
Rwpos38_91 in38 sp91 11140.846016
Rwpos38_92 in38 sp92 3183.098862
Rwpos38_93 in38 sp93 3183.098862
Rwpos38_94 in38 sp94 3183.098862
Rwpos38_95 in38 sp95 11140.846016
Rwpos38_96 in38 sp96 11140.846016
Rwpos38_97 in38 sp97 11140.846016
Rwpos38_98 in38 sp98 3183.098862
Rwpos38_99 in38 sp99 3183.098862
Rwpos38_100 in38 sp100 3183.098862
Rwpos39_1 in39 sp1 11140.846016
Rwpos39_2 in39 sp2 3183.098862
Rwpos39_3 in39 sp3 11140.846016
Rwpos39_4 in39 sp4 3183.098862
Rwpos39_5 in39 sp5 3183.098862
Rwpos39_6 in39 sp6 3183.098862
Rwpos39_7 in39 sp7 3183.098862
Rwpos39_8 in39 sp8 11140.846016
Rwpos39_9 in39 sp9 3183.098862
Rwpos39_10 in39 sp10 3183.098862
Rwpos39_11 in39 sp11 11140.846016
Rwpos39_12 in39 sp12 3183.098862
Rwpos39_13 in39 sp13 3183.098862
Rwpos39_14 in39 sp14 3183.098862
Rwpos39_15 in39 sp15 11140.846016
Rwpos39_16 in39 sp16 3183.098862
Rwpos39_17 in39 sp17 3183.098862
Rwpos39_18 in39 sp18 3183.098862
Rwpos39_19 in39 sp19 3183.098862
Rwpos39_20 in39 sp20 11140.846016
Rwpos39_21 in39 sp21 3183.098862
Rwpos39_22 in39 sp22 3183.098862
Rwpos39_23 in39 sp23 11140.846016
Rwpos39_24 in39 sp24 3183.098862
Rwpos39_25 in39 sp25 11140.846016
Rwpos39_26 in39 sp26 3183.098862
Rwpos39_27 in39 sp27 11140.846016
Rwpos39_28 in39 sp28 11140.846016
Rwpos39_29 in39 sp29 11140.846016
Rwpos39_30 in39 sp30 3183.098862
Rwpos39_31 in39 sp31 3183.098862
Rwpos39_32 in39 sp32 3183.098862
Rwpos39_33 in39 sp33 3183.098862
Rwpos39_34 in39 sp34 3183.098862
Rwpos39_35 in39 sp35 11140.846016
Rwpos39_36 in39 sp36 11140.846016
Rwpos39_37 in39 sp37 3183.098862
Rwpos39_38 in39 sp38 11140.846016
Rwpos39_39 in39 sp39 3183.098862
Rwpos39_40 in39 sp40 3183.098862
Rwpos39_41 in39 sp41 3183.098862
Rwpos39_42 in39 sp42 3183.098862
Rwpos39_43 in39 sp43 11140.846016
Rwpos39_44 in39 sp44 11140.846016
Rwpos39_45 in39 sp45 11140.846016
Rwpos39_46 in39 sp46 3183.098862
Rwpos39_47 in39 sp47 3183.098862
Rwpos39_48 in39 sp48 11140.846016
Rwpos39_49 in39 sp49 11140.846016
Rwpos39_50 in39 sp50 3183.098862
Rwpos39_51 in39 sp51 11140.846016
Rwpos39_52 in39 sp52 11140.846016
Rwpos39_53 in39 sp53 3183.098862
Rwpos39_54 in39 sp54 3183.098862
Rwpos39_55 in39 sp55 11140.846016
Rwpos39_56 in39 sp56 3183.098862
Rwpos39_57 in39 sp57 11140.846016
Rwpos39_58 in39 sp58 3183.098862
Rwpos39_59 in39 sp59 11140.846016
Rwpos39_60 in39 sp60 11140.846016
Rwpos39_61 in39 sp61 3183.098862
Rwpos39_62 in39 sp62 3183.098862
Rwpos39_63 in39 sp63 3183.098862
Rwpos39_64 in39 sp64 3183.098862
Rwpos39_65 in39 sp65 11140.846016
Rwpos39_66 in39 sp66 3183.098862
Rwpos39_67 in39 sp67 3183.098862
Rwpos39_68 in39 sp68 11140.846016
Rwpos39_69 in39 sp69 3183.098862
Rwpos39_70 in39 sp70 3183.098862
Rwpos39_71 in39 sp71 11140.846016
Rwpos39_72 in39 sp72 3183.098862
Rwpos39_73 in39 sp73 11140.846016
Rwpos39_74 in39 sp74 3183.098862
Rwpos39_75 in39 sp75 3183.098862
Rwpos39_76 in39 sp76 3183.098862
Rwpos39_77 in39 sp77 11140.846016
Rwpos39_78 in39 sp78 3183.098862
Rwpos39_79 in39 sp79 3183.098862
Rwpos39_80 in39 sp80 3183.098862
Rwpos39_81 in39 sp81 11140.846016
Rwpos39_82 in39 sp82 3183.098862
Rwpos39_83 in39 sp83 11140.846016
Rwpos39_84 in39 sp84 3183.098862
Rwpos39_85 in39 sp85 11140.846016
Rwpos39_86 in39 sp86 11140.846016
Rwpos39_87 in39 sp87 11140.846016
Rwpos39_88 in39 sp88 3183.098862
Rwpos39_89 in39 sp89 11140.846016
Rwpos39_90 in39 sp90 3183.098862
Rwpos39_91 in39 sp91 3183.098862
Rwpos39_92 in39 sp92 11140.846016
Rwpos39_93 in39 sp93 3183.098862
Rwpos39_94 in39 sp94 3183.098862
Rwpos39_95 in39 sp95 11140.846016
Rwpos39_96 in39 sp96 3183.098862
Rwpos39_97 in39 sp97 3183.098862
Rwpos39_98 in39 sp98 3183.098862
Rwpos39_99 in39 sp99 3183.098862
Rwpos39_100 in39 sp100 3183.098862
Rwpos40_1 in40 sp1 11140.846016
Rwpos40_2 in40 sp2 3183.098862
Rwpos40_3 in40 sp3 3183.098862
Rwpos40_4 in40 sp4 3183.098862
Rwpos40_5 in40 sp5 11140.846016
Rwpos40_6 in40 sp6 11140.846016
Rwpos40_7 in40 sp7 3183.098862
Rwpos40_8 in40 sp8 3183.098862
Rwpos40_9 in40 sp9 11140.846016
Rwpos40_10 in40 sp10 3183.098862
Rwpos40_11 in40 sp11 3183.098862
Rwpos40_12 in40 sp12 11140.846016
Rwpos40_13 in40 sp13 3183.098862
Rwpos40_14 in40 sp14 3183.098862
Rwpos40_15 in40 sp15 11140.846016
Rwpos40_16 in40 sp16 3183.098862
Rwpos40_17 in40 sp17 11140.846016
Rwpos40_18 in40 sp18 11140.846016
Rwpos40_19 in40 sp19 3183.098862
Rwpos40_20 in40 sp20 3183.098862
Rwpos40_21 in40 sp21 11140.846016
Rwpos40_22 in40 sp22 3183.098862
Rwpos40_23 in40 sp23 3183.098862
Rwpos40_24 in40 sp24 11140.846016
Rwpos40_25 in40 sp25 3183.098862
Rwpos40_26 in40 sp26 3183.098862
Rwpos40_27 in40 sp27 3183.098862
Rwpos40_28 in40 sp28 3183.098862
Rwpos40_29 in40 sp29 11140.846016
Rwpos40_30 in40 sp30 3183.098862
Rwpos40_31 in40 sp31 11140.846016
Rwpos40_32 in40 sp32 11140.846016
Rwpos40_33 in40 sp33 11140.846016
Rwpos40_34 in40 sp34 3183.098862
Rwpos40_35 in40 sp35 11140.846016
Rwpos40_36 in40 sp36 3183.098862
Rwpos40_37 in40 sp37 11140.846016
Rwpos40_38 in40 sp38 11140.846016
Rwpos40_39 in40 sp39 3183.098862
Rwpos40_40 in40 sp40 3183.098862
Rwpos40_41 in40 sp41 3183.098862
Rwpos40_42 in40 sp42 3183.098862
Rwpos40_43 in40 sp43 11140.846016
Rwpos40_44 in40 sp44 3183.098862
Rwpos40_45 in40 sp45 11140.846016
Rwpos40_46 in40 sp46 3183.098862
Rwpos40_47 in40 sp47 3183.098862
Rwpos40_48 in40 sp48 3183.098862
Rwpos40_49 in40 sp49 11140.846016
Rwpos40_50 in40 sp50 3183.098862
Rwpos40_51 in40 sp51 3183.098862
Rwpos40_52 in40 sp52 3183.098862
Rwpos40_53 in40 sp53 11140.846016
Rwpos40_54 in40 sp54 11140.846016
Rwpos40_55 in40 sp55 3183.098862
Rwpos40_56 in40 sp56 3183.098862
Rwpos40_57 in40 sp57 3183.098862
Rwpos40_58 in40 sp58 3183.098862
Rwpos40_59 in40 sp59 11140.846016
Rwpos40_60 in40 sp60 3183.098862
Rwpos40_61 in40 sp61 11140.846016
Rwpos40_62 in40 sp62 3183.098862
Rwpos40_63 in40 sp63 3183.098862
Rwpos40_64 in40 sp64 3183.098862
Rwpos40_65 in40 sp65 11140.846016
Rwpos40_66 in40 sp66 11140.846016
Rwpos40_67 in40 sp67 3183.098862
Rwpos40_68 in40 sp68 3183.098862
Rwpos40_69 in40 sp69 3183.098862
Rwpos40_70 in40 sp70 3183.098862
Rwpos40_71 in40 sp71 11140.846016
Rwpos40_72 in40 sp72 3183.098862
Rwpos40_73 in40 sp73 11140.846016
Rwpos40_74 in40 sp74 11140.846016
Rwpos40_75 in40 sp75 11140.846016
Rwpos40_76 in40 sp76 3183.098862
Rwpos40_77 in40 sp77 11140.846016
Rwpos40_78 in40 sp78 3183.098862
Rwpos40_79 in40 sp79 3183.098862
Rwpos40_80 in40 sp80 3183.098862
Rwpos40_81 in40 sp81 11140.846016
Rwpos40_82 in40 sp82 3183.098862
Rwpos40_83 in40 sp83 3183.098862
Rwpos40_84 in40 sp84 3183.098862
Rwpos40_85 in40 sp85 3183.098862
Rwpos40_86 in40 sp86 3183.098862
Rwpos40_87 in40 sp87 3183.098862
Rwpos40_88 in40 sp88 11140.846016
Rwpos40_89 in40 sp89 3183.098862
Rwpos40_90 in40 sp90 3183.098862
Rwpos40_91 in40 sp91 11140.846016
Rwpos40_92 in40 sp92 11140.846016
Rwpos40_93 in40 sp93 11140.846016
Rwpos40_94 in40 sp94 3183.098862
Rwpos40_95 in40 sp95 3183.098862
Rwpos40_96 in40 sp96 3183.098862
Rwpos40_97 in40 sp97 11140.846016
Rwpos40_98 in40 sp98 3183.098862
Rwpos40_99 in40 sp99 3183.098862
Rwpos40_100 in40 sp100 3183.098862
Rwpos41_1 in41 sp1 11140.846016
Rwpos41_2 in41 sp2 3183.098862
Rwpos41_3 in41 sp3 3183.098862
Rwpos41_4 in41 sp4 11140.846016
Rwpos41_5 in41 sp5 3183.098862
Rwpos41_6 in41 sp6 3183.098862
Rwpos41_7 in41 sp7 11140.846016
Rwpos41_8 in41 sp8 3183.098862
Rwpos41_9 in41 sp9 11140.846016
Rwpos41_10 in41 sp10 11140.846016
Rwpos41_11 in41 sp11 3183.098862
Rwpos41_12 in41 sp12 3183.098862
Rwpos41_13 in41 sp13 11140.846016
Rwpos41_14 in41 sp14 3183.098862
Rwpos41_15 in41 sp15 3183.098862
Rwpos41_16 in41 sp16 11140.846016
Rwpos41_17 in41 sp17 11140.846016
Rwpos41_18 in41 sp18 11140.846016
Rwpos41_19 in41 sp19 3183.098862
Rwpos41_20 in41 sp20 11140.846016
Rwpos41_21 in41 sp21 3183.098862
Rwpos41_22 in41 sp22 3183.098862
Rwpos41_23 in41 sp23 3183.098862
Rwpos41_24 in41 sp24 11140.846016
Rwpos41_25 in41 sp25 3183.098862
Rwpos41_26 in41 sp26 11140.846016
Rwpos41_27 in41 sp27 11140.846016
Rwpos41_28 in41 sp28 3183.098862
Rwpos41_29 in41 sp29 3183.098862
Rwpos41_30 in41 sp30 11140.846016
Rwpos41_31 in41 sp31 3183.098862
Rwpos41_32 in41 sp32 11140.846016
Rwpos41_33 in41 sp33 3183.098862
Rwpos41_34 in41 sp34 3183.098862
Rwpos41_35 in41 sp35 11140.846016
Rwpos41_36 in41 sp36 3183.098862
Rwpos41_37 in41 sp37 3183.098862
Rwpos41_38 in41 sp38 3183.098862
Rwpos41_39 in41 sp39 3183.098862
Rwpos41_40 in41 sp40 3183.098862
Rwpos41_41 in41 sp41 3183.098862
Rwpos41_42 in41 sp42 3183.098862
Rwpos41_43 in41 sp43 11140.846016
Rwpos41_44 in41 sp44 3183.098862
Rwpos41_45 in41 sp45 3183.098862
Rwpos41_46 in41 sp46 11140.846016
Rwpos41_47 in41 sp47 3183.098862
Rwpos41_48 in41 sp48 3183.098862
Rwpos41_49 in41 sp49 11140.846016
Rwpos41_50 in41 sp50 11140.846016
Rwpos41_51 in41 sp51 11140.846016
Rwpos41_52 in41 sp52 11140.846016
Rwpos41_53 in41 sp53 11140.846016
Rwpos41_54 in41 sp54 3183.098862
Rwpos41_55 in41 sp55 3183.098862
Rwpos41_56 in41 sp56 11140.846016
Rwpos41_57 in41 sp57 11140.846016
Rwpos41_58 in41 sp58 11140.846016
Rwpos41_59 in41 sp59 11140.846016
Rwpos41_60 in41 sp60 3183.098862
Rwpos41_61 in41 sp61 11140.846016
Rwpos41_62 in41 sp62 11140.846016
Rwpos41_63 in41 sp63 3183.098862
Rwpos41_64 in41 sp64 3183.098862
Rwpos41_65 in41 sp65 11140.846016
Rwpos41_66 in41 sp66 3183.098862
Rwpos41_67 in41 sp67 3183.098862
Rwpos41_68 in41 sp68 11140.846016
Rwpos41_69 in41 sp69 11140.846016
Rwpos41_70 in41 sp70 3183.098862
Rwpos41_71 in41 sp71 3183.098862
Rwpos41_72 in41 sp72 3183.098862
Rwpos41_73 in41 sp73 11140.846016
Rwpos41_74 in41 sp74 11140.846016
Rwpos41_75 in41 sp75 11140.846016
Rwpos41_76 in41 sp76 3183.098862
Rwpos41_77 in41 sp77 11140.846016
Rwpos41_78 in41 sp78 11140.846016
Rwpos41_79 in41 sp79 11140.846016
Rwpos41_80 in41 sp80 11140.846016
Rwpos41_81 in41 sp81 11140.846016
Rwpos41_82 in41 sp82 3183.098862
Rwpos41_83 in41 sp83 11140.846016
Rwpos41_84 in41 sp84 11140.846016
Rwpos41_85 in41 sp85 3183.098862
Rwpos41_86 in41 sp86 3183.098862
Rwpos41_87 in41 sp87 3183.098862
Rwpos41_88 in41 sp88 11140.846016
Rwpos41_89 in41 sp89 3183.098862
Rwpos41_90 in41 sp90 3183.098862
Rwpos41_91 in41 sp91 11140.846016
Rwpos41_92 in41 sp92 3183.098862
Rwpos41_93 in41 sp93 3183.098862
Rwpos41_94 in41 sp94 3183.098862
Rwpos41_95 in41 sp95 11140.846016
Rwpos41_96 in41 sp96 3183.098862
Rwpos41_97 in41 sp97 11140.846016
Rwpos41_98 in41 sp98 3183.098862
Rwpos41_99 in41 sp99 3183.098862
Rwpos41_100 in41 sp100 11140.846016
Rwpos42_1 in42 sp1 3183.098862
Rwpos42_2 in42 sp2 3183.098862
Rwpos42_3 in42 sp3 11140.846016
Rwpos42_4 in42 sp4 3183.098862
Rwpos42_5 in42 sp5 3183.098862
Rwpos42_6 in42 sp6 11140.846016
Rwpos42_7 in42 sp7 11140.846016
Rwpos42_8 in42 sp8 3183.098862
Rwpos42_9 in42 sp9 3183.098862
Rwpos42_10 in42 sp10 3183.098862
Rwpos42_11 in42 sp11 11140.846016
Rwpos42_12 in42 sp12 11140.846016
Rwpos42_13 in42 sp13 11140.846016
Rwpos42_14 in42 sp14 11140.846016
Rwpos42_15 in42 sp15 3183.098862
Rwpos42_16 in42 sp16 11140.846016
Rwpos42_17 in42 sp17 11140.846016
Rwpos42_18 in42 sp18 3183.098862
Rwpos42_19 in42 sp19 3183.098862
Rwpos42_20 in42 sp20 3183.098862
Rwpos42_21 in42 sp21 11140.846016
Rwpos42_22 in42 sp22 11140.846016
Rwpos42_23 in42 sp23 11140.846016
Rwpos42_24 in42 sp24 3183.098862
Rwpos42_25 in42 sp25 11140.846016
Rwpos42_26 in42 sp26 11140.846016
Rwpos42_27 in42 sp27 11140.846016
Rwpos42_28 in42 sp28 11140.846016
Rwpos42_29 in42 sp29 11140.846016
Rwpos42_30 in42 sp30 3183.098862
Rwpos42_31 in42 sp31 3183.098862
Rwpos42_32 in42 sp32 3183.098862
Rwpos42_33 in42 sp33 11140.846016
Rwpos42_34 in42 sp34 11140.846016
Rwpos42_35 in42 sp35 3183.098862
Rwpos42_36 in42 sp36 3183.098862
Rwpos42_37 in42 sp37 3183.098862
Rwpos42_38 in42 sp38 3183.098862
Rwpos42_39 in42 sp39 3183.098862
Rwpos42_40 in42 sp40 3183.098862
Rwpos42_41 in42 sp41 3183.098862
Rwpos42_42 in42 sp42 3183.098862
Rwpos42_43 in42 sp43 11140.846016
Rwpos42_44 in42 sp44 11140.846016
Rwpos42_45 in42 sp45 3183.098862
Rwpos42_46 in42 sp46 11140.846016
Rwpos42_47 in42 sp47 3183.098862
Rwpos42_48 in42 sp48 11140.846016
Rwpos42_49 in42 sp49 11140.846016
Rwpos42_50 in42 sp50 3183.098862
Rwpos42_51 in42 sp51 3183.098862
Rwpos42_52 in42 sp52 3183.098862
Rwpos42_53 in42 sp53 11140.846016
Rwpos42_54 in42 sp54 3183.098862
Rwpos42_55 in42 sp55 3183.098862
Rwpos42_56 in42 sp56 3183.098862
Rwpos42_57 in42 sp57 11140.846016
Rwpos42_58 in42 sp58 11140.846016
Rwpos42_59 in42 sp59 11140.846016
Rwpos42_60 in42 sp60 3183.098862
Rwpos42_61 in42 sp61 3183.098862
Rwpos42_62 in42 sp62 11140.846016
Rwpos42_63 in42 sp63 11140.846016
Rwpos42_64 in42 sp64 11140.846016
Rwpos42_65 in42 sp65 11140.846016
Rwpos42_66 in42 sp66 11140.846016
Rwpos42_67 in42 sp67 3183.098862
Rwpos42_68 in42 sp68 3183.098862
Rwpos42_69 in42 sp69 11140.846016
Rwpos42_70 in42 sp70 3183.098862
Rwpos42_71 in42 sp71 3183.098862
Rwpos42_72 in42 sp72 3183.098862
Rwpos42_73 in42 sp73 11140.846016
Rwpos42_74 in42 sp74 3183.098862
Rwpos42_75 in42 sp75 11140.846016
Rwpos42_76 in42 sp76 3183.098862
Rwpos42_77 in42 sp77 3183.098862
Rwpos42_78 in42 sp78 3183.098862
Rwpos42_79 in42 sp79 3183.098862
Rwpos42_80 in42 sp80 3183.098862
Rwpos42_81 in42 sp81 11140.846016
Rwpos42_82 in42 sp82 3183.098862
Rwpos42_83 in42 sp83 3183.098862
Rwpos42_84 in42 sp84 11140.846016
Rwpos42_85 in42 sp85 11140.846016
Rwpos42_86 in42 sp86 3183.098862
Rwpos42_87 in42 sp87 3183.098862
Rwpos42_88 in42 sp88 3183.098862
Rwpos42_89 in42 sp89 11140.846016
Rwpos42_90 in42 sp90 11140.846016
Rwpos42_91 in42 sp91 11140.846016
Rwpos42_92 in42 sp92 3183.098862
Rwpos42_93 in42 sp93 3183.098862
Rwpos42_94 in42 sp94 11140.846016
Rwpos42_95 in42 sp95 3183.098862
Rwpos42_96 in42 sp96 3183.098862
Rwpos42_97 in42 sp97 11140.846016
Rwpos42_98 in42 sp98 3183.098862
Rwpos42_99 in42 sp99 3183.098862
Rwpos42_100 in42 sp100 3183.098862
Rwpos43_1 in43 sp1 3183.098862
Rwpos43_2 in43 sp2 3183.098862
Rwpos43_3 in43 sp3 3183.098862
Rwpos43_4 in43 sp4 3183.098862
Rwpos43_5 in43 sp5 11140.846016
Rwpos43_6 in43 sp6 11140.846016
Rwpos43_7 in43 sp7 3183.098862
Rwpos43_8 in43 sp8 11140.846016
Rwpos43_9 in43 sp9 3183.098862
Rwpos43_10 in43 sp10 3183.098862
Rwpos43_11 in43 sp11 3183.098862
Rwpos43_12 in43 sp12 11140.846016
Rwpos43_13 in43 sp13 11140.846016
Rwpos43_14 in43 sp14 3183.098862
Rwpos43_15 in43 sp15 3183.098862
Rwpos43_16 in43 sp16 11140.846016
Rwpos43_17 in43 sp17 11140.846016
Rwpos43_18 in43 sp18 3183.098862
Rwpos43_19 in43 sp19 3183.098862
Rwpos43_20 in43 sp20 11140.846016
Rwpos43_21 in43 sp21 11140.846016
Rwpos43_22 in43 sp22 11140.846016
Rwpos43_23 in43 sp23 11140.846016
Rwpos43_24 in43 sp24 11140.846016
Rwpos43_25 in43 sp25 3183.098862
Rwpos43_26 in43 sp26 3183.098862
Rwpos43_27 in43 sp27 3183.098862
Rwpos43_28 in43 sp28 3183.098862
Rwpos43_29 in43 sp29 11140.846016
Rwpos43_30 in43 sp30 3183.098862
Rwpos43_31 in43 sp31 3183.098862
Rwpos43_32 in43 sp32 11140.846016
Rwpos43_33 in43 sp33 11140.846016
Rwpos43_34 in43 sp34 3183.098862
Rwpos43_35 in43 sp35 3183.098862
Rwpos43_36 in43 sp36 3183.098862
Rwpos43_37 in43 sp37 11140.846016
Rwpos43_38 in43 sp38 11140.846016
Rwpos43_39 in43 sp39 11140.846016
Rwpos43_40 in43 sp40 3183.098862
Rwpos43_41 in43 sp41 11140.846016
Rwpos43_42 in43 sp42 3183.098862
Rwpos43_43 in43 sp43 11140.846016
Rwpos43_44 in43 sp44 11140.846016
Rwpos43_45 in43 sp45 11140.846016
Rwpos43_46 in43 sp46 3183.098862
Rwpos43_47 in43 sp47 11140.846016
Rwpos43_48 in43 sp48 3183.098862
Rwpos43_49 in43 sp49 3183.098862
Rwpos43_50 in43 sp50 3183.098862
Rwpos43_51 in43 sp51 3183.098862
Rwpos43_52 in43 sp52 11140.846016
Rwpos43_53 in43 sp53 11140.846016
Rwpos43_54 in43 sp54 11140.846016
Rwpos43_55 in43 sp55 11140.846016
Rwpos43_56 in43 sp56 11140.846016
Rwpos43_57 in43 sp57 11140.846016
Rwpos43_58 in43 sp58 3183.098862
Rwpos43_59 in43 sp59 11140.846016
Rwpos43_60 in43 sp60 11140.846016
Rwpos43_61 in43 sp61 3183.098862
Rwpos43_62 in43 sp62 3183.098862
Rwpos43_63 in43 sp63 11140.846016
Rwpos43_64 in43 sp64 11140.846016
Rwpos43_65 in43 sp65 11140.846016
Rwpos43_66 in43 sp66 3183.098862
Rwpos43_67 in43 sp67 11140.846016
Rwpos43_68 in43 sp68 11140.846016
Rwpos43_69 in43 sp69 3183.098862
Rwpos43_70 in43 sp70 11140.846016
Rwpos43_71 in43 sp71 11140.846016
Rwpos43_72 in43 sp72 3183.098862
Rwpos43_73 in43 sp73 11140.846016
Rwpos43_74 in43 sp74 3183.098862
Rwpos43_75 in43 sp75 11140.846016
Rwpos43_76 in43 sp76 11140.846016
Rwpos43_77 in43 sp77 11140.846016
Rwpos43_78 in43 sp78 3183.098862
Rwpos43_79 in43 sp79 11140.846016
Rwpos43_80 in43 sp80 3183.098862
Rwpos43_81 in43 sp81 3183.098862
Rwpos43_82 in43 sp82 3183.098862
Rwpos43_83 in43 sp83 11140.846016
Rwpos43_84 in43 sp84 11140.846016
Rwpos43_85 in43 sp85 3183.098862
Rwpos43_86 in43 sp86 3183.098862
Rwpos43_87 in43 sp87 11140.846016
Rwpos43_88 in43 sp88 3183.098862
Rwpos43_89 in43 sp89 11140.846016
Rwpos43_90 in43 sp90 3183.098862
Rwpos43_91 in43 sp91 3183.098862
Rwpos43_92 in43 sp92 11140.846016
Rwpos43_93 in43 sp93 11140.846016
Rwpos43_94 in43 sp94 3183.098862
Rwpos43_95 in43 sp95 11140.846016
Rwpos43_96 in43 sp96 11140.846016
Rwpos43_97 in43 sp97 3183.098862
Rwpos43_98 in43 sp98 3183.098862
Rwpos43_99 in43 sp99 11140.846016
Rwpos43_100 in43 sp100 11140.846016
Rwpos44_1 in44 sp1 3183.098862
Rwpos44_2 in44 sp2 3183.098862
Rwpos44_3 in44 sp3 11140.846016
Rwpos44_4 in44 sp4 3183.098862
Rwpos44_5 in44 sp5 11140.846016
Rwpos44_6 in44 sp6 3183.098862
Rwpos44_7 in44 sp7 3183.098862
Rwpos44_8 in44 sp8 11140.846016
Rwpos44_9 in44 sp9 11140.846016
Rwpos44_10 in44 sp10 3183.098862
Rwpos44_11 in44 sp11 11140.846016
Rwpos44_12 in44 sp12 11140.846016
Rwpos44_13 in44 sp13 3183.098862
Rwpos44_14 in44 sp14 3183.098862
Rwpos44_15 in44 sp15 3183.098862
Rwpos44_16 in44 sp16 11140.846016
Rwpos44_17 in44 sp17 3183.098862
Rwpos44_18 in44 sp18 3183.098862
Rwpos44_19 in44 sp19 11140.846016
Rwpos44_20 in44 sp20 3183.098862
Rwpos44_21 in44 sp21 11140.846016
Rwpos44_22 in44 sp22 3183.098862
Rwpos44_23 in44 sp23 3183.098862
Rwpos44_24 in44 sp24 11140.846016
Rwpos44_25 in44 sp25 11140.846016
Rwpos44_26 in44 sp26 3183.098862
Rwpos44_27 in44 sp27 11140.846016
Rwpos44_28 in44 sp28 11140.846016
Rwpos44_29 in44 sp29 11140.846016
Rwpos44_30 in44 sp30 3183.098862
Rwpos44_31 in44 sp31 11140.846016
Rwpos44_32 in44 sp32 11140.846016
Rwpos44_33 in44 sp33 3183.098862
Rwpos44_34 in44 sp34 3183.098862
Rwpos44_35 in44 sp35 11140.846016
Rwpos44_36 in44 sp36 3183.098862
Rwpos44_37 in44 sp37 11140.846016
Rwpos44_38 in44 sp38 11140.846016
Rwpos44_39 in44 sp39 11140.846016
Rwpos44_40 in44 sp40 3183.098862
Rwpos44_41 in44 sp41 11140.846016
Rwpos44_42 in44 sp42 3183.098862
Rwpos44_43 in44 sp43 3183.098862
Rwpos44_44 in44 sp44 11140.846016
Rwpos44_45 in44 sp45 11140.846016
Rwpos44_46 in44 sp46 3183.098862
Rwpos44_47 in44 sp47 11140.846016
Rwpos44_48 in44 sp48 11140.846016
Rwpos44_49 in44 sp49 3183.098862
Rwpos44_50 in44 sp50 11140.846016
Rwpos44_51 in44 sp51 11140.846016
Rwpos44_52 in44 sp52 3183.098862
Rwpos44_53 in44 sp53 11140.846016
Rwpos44_54 in44 sp54 11140.846016
Rwpos44_55 in44 sp55 3183.098862
Rwpos44_56 in44 sp56 11140.846016
Rwpos44_57 in44 sp57 3183.098862
Rwpos44_58 in44 sp58 3183.098862
Rwpos44_59 in44 sp59 11140.846016
Rwpos44_60 in44 sp60 3183.098862
Rwpos44_61 in44 sp61 3183.098862
Rwpos44_62 in44 sp62 3183.098862
Rwpos44_63 in44 sp63 3183.098862
Rwpos44_64 in44 sp64 11140.846016
Rwpos44_65 in44 sp65 3183.098862
Rwpos44_66 in44 sp66 11140.846016
Rwpos44_67 in44 sp67 11140.846016
Rwpos44_68 in44 sp68 3183.098862
Rwpos44_69 in44 sp69 11140.846016
Rwpos44_70 in44 sp70 11140.846016
Rwpos44_71 in44 sp71 3183.098862
Rwpos44_72 in44 sp72 3183.098862
Rwpos44_73 in44 sp73 3183.098862
Rwpos44_74 in44 sp74 3183.098862
Rwpos44_75 in44 sp75 11140.846016
Rwpos44_76 in44 sp76 3183.098862
Rwpos44_77 in44 sp77 11140.846016
Rwpos44_78 in44 sp78 3183.098862
Rwpos44_79 in44 sp79 11140.846016
Rwpos44_80 in44 sp80 11140.846016
Rwpos44_81 in44 sp81 11140.846016
Rwpos44_82 in44 sp82 3183.098862
Rwpos44_83 in44 sp83 3183.098862
Rwpos44_84 in44 sp84 3183.098862
Rwpos44_85 in44 sp85 11140.846016
Rwpos44_86 in44 sp86 11140.846016
Rwpos44_87 in44 sp87 3183.098862
Rwpos44_88 in44 sp88 3183.098862
Rwpos44_89 in44 sp89 11140.846016
Rwpos44_90 in44 sp90 3183.098862
Rwpos44_91 in44 sp91 3183.098862
Rwpos44_92 in44 sp92 11140.846016
Rwpos44_93 in44 sp93 11140.846016
Rwpos44_94 in44 sp94 3183.098862
Rwpos44_95 in44 sp95 3183.098862
Rwpos44_96 in44 sp96 11140.846016
Rwpos44_97 in44 sp97 11140.846016
Rwpos44_98 in44 sp98 11140.846016
Rwpos44_99 in44 sp99 11140.846016
Rwpos44_100 in44 sp100 3183.098862
Rwpos45_1 in45 sp1 3183.098862
Rwpos45_2 in45 sp2 11140.846016
Rwpos45_3 in45 sp3 3183.098862
Rwpos45_4 in45 sp4 3183.098862
Rwpos45_5 in45 sp5 3183.098862
Rwpos45_6 in45 sp6 3183.098862
Rwpos45_7 in45 sp7 11140.846016
Rwpos45_8 in45 sp8 3183.098862
Rwpos45_9 in45 sp9 11140.846016
Rwpos45_10 in45 sp10 3183.098862
Rwpos45_11 in45 sp11 3183.098862
Rwpos45_12 in45 sp12 3183.098862
Rwpos45_13 in45 sp13 11140.846016
Rwpos45_14 in45 sp14 11140.846016
Rwpos45_15 in45 sp15 11140.846016
Rwpos45_16 in45 sp16 3183.098862
Rwpos45_17 in45 sp17 3183.098862
Rwpos45_18 in45 sp18 11140.846016
Rwpos45_19 in45 sp19 3183.098862
Rwpos45_20 in45 sp20 3183.098862
Rwpos45_21 in45 sp21 11140.846016
Rwpos45_22 in45 sp22 3183.098862
Rwpos45_23 in45 sp23 11140.846016
Rwpos45_24 in45 sp24 3183.098862
Rwpos45_25 in45 sp25 11140.846016
Rwpos45_26 in45 sp26 3183.098862
Rwpos45_27 in45 sp27 3183.098862
Rwpos45_28 in45 sp28 3183.098862
Rwpos45_29 in45 sp29 11140.846016
Rwpos45_30 in45 sp30 3183.098862
Rwpos45_31 in45 sp31 3183.098862
Rwpos45_32 in45 sp32 3183.098862
Rwpos45_33 in45 sp33 3183.098862
Rwpos45_34 in45 sp34 3183.098862
Rwpos45_35 in45 sp35 3183.098862
Rwpos45_36 in45 sp36 3183.098862
Rwpos45_37 in45 sp37 3183.098862
Rwpos45_38 in45 sp38 3183.098862
Rwpos45_39 in45 sp39 11140.846016
Rwpos45_40 in45 sp40 11140.846016
Rwpos45_41 in45 sp41 11140.846016
Rwpos45_42 in45 sp42 3183.098862
Rwpos45_43 in45 sp43 11140.846016
Rwpos45_44 in45 sp44 11140.846016
Rwpos45_45 in45 sp45 11140.846016
Rwpos45_46 in45 sp46 3183.098862
Rwpos45_47 in45 sp47 3183.098862
Rwpos45_48 in45 sp48 3183.098862
Rwpos45_49 in45 sp49 11140.846016
Rwpos45_50 in45 sp50 11140.846016
Rwpos45_51 in45 sp51 11140.846016
Rwpos45_52 in45 sp52 11140.846016
Rwpos45_53 in45 sp53 11140.846016
Rwpos45_54 in45 sp54 11140.846016
Rwpos45_55 in45 sp55 11140.846016
Rwpos45_56 in45 sp56 3183.098862
Rwpos45_57 in45 sp57 3183.098862
Rwpos45_58 in45 sp58 3183.098862
Rwpos45_59 in45 sp59 11140.846016
Rwpos45_60 in45 sp60 3183.098862
Rwpos45_61 in45 sp61 3183.098862
Rwpos45_62 in45 sp62 11140.846016
Rwpos45_63 in45 sp63 3183.098862
Rwpos45_64 in45 sp64 3183.098862
Rwpos45_65 in45 sp65 3183.098862
Rwpos45_66 in45 sp66 11140.846016
Rwpos45_67 in45 sp67 3183.098862
Rwpos45_68 in45 sp68 11140.846016
Rwpos45_69 in45 sp69 11140.846016
Rwpos45_70 in45 sp70 3183.098862
Rwpos45_71 in45 sp71 3183.098862
Rwpos45_72 in45 sp72 3183.098862
Rwpos45_73 in45 sp73 3183.098862
Rwpos45_74 in45 sp74 3183.098862
Rwpos45_75 in45 sp75 3183.098862
Rwpos45_76 in45 sp76 11140.846016
Rwpos45_77 in45 sp77 11140.846016
Rwpos45_78 in45 sp78 11140.846016
Rwpos45_79 in45 sp79 3183.098862
Rwpos45_80 in45 sp80 11140.846016
Rwpos45_81 in45 sp81 3183.098862
Rwpos45_82 in45 sp82 3183.098862
Rwpos45_83 in45 sp83 11140.846016
Rwpos45_84 in45 sp84 11140.846016
Rwpos45_85 in45 sp85 3183.098862
Rwpos45_86 in45 sp86 11140.846016
Rwpos45_87 in45 sp87 3183.098862
Rwpos45_88 in45 sp88 3183.098862
Rwpos45_89 in45 sp89 3183.098862
Rwpos45_90 in45 sp90 3183.098862
Rwpos45_91 in45 sp91 11140.846016
Rwpos45_92 in45 sp92 3183.098862
Rwpos45_93 in45 sp93 11140.846016
Rwpos45_94 in45 sp94 11140.846016
Rwpos45_95 in45 sp95 3183.098862
Rwpos45_96 in45 sp96 3183.098862
Rwpos45_97 in45 sp97 11140.846016
Rwpos45_98 in45 sp98 3183.098862
Rwpos45_99 in45 sp99 3183.098862
Rwpos45_100 in45 sp100 3183.098862
Rwpos46_1 in46 sp1 11140.846016
Rwpos46_2 in46 sp2 3183.098862
Rwpos46_3 in46 sp3 11140.846016
Rwpos46_4 in46 sp4 3183.098862
Rwpos46_5 in46 sp5 3183.098862
Rwpos46_6 in46 sp6 11140.846016
Rwpos46_7 in46 sp7 3183.098862
Rwpos46_8 in46 sp8 11140.846016
Rwpos46_9 in46 sp9 11140.846016
Rwpos46_10 in46 sp10 11140.846016
Rwpos46_11 in46 sp11 11140.846016
Rwpos46_12 in46 sp12 11140.846016
Rwpos46_13 in46 sp13 11140.846016
Rwpos46_14 in46 sp14 3183.098862
Rwpos46_15 in46 sp15 3183.098862
Rwpos46_16 in46 sp16 11140.846016
Rwpos46_17 in46 sp17 3183.098862
Rwpos46_18 in46 sp18 11140.846016
Rwpos46_19 in46 sp19 3183.098862
Rwpos46_20 in46 sp20 11140.846016
Rwpos46_21 in46 sp21 11140.846016
Rwpos46_22 in46 sp22 3183.098862
Rwpos46_23 in46 sp23 3183.098862
Rwpos46_24 in46 sp24 11140.846016
Rwpos46_25 in46 sp25 11140.846016
Rwpos46_26 in46 sp26 3183.098862
Rwpos46_27 in46 sp27 11140.846016
Rwpos46_28 in46 sp28 11140.846016
Rwpos46_29 in46 sp29 3183.098862
Rwpos46_30 in46 sp30 3183.098862
Rwpos46_31 in46 sp31 11140.846016
Rwpos46_32 in46 sp32 3183.098862
Rwpos46_33 in46 sp33 3183.098862
Rwpos46_34 in46 sp34 11140.846016
Rwpos46_35 in46 sp35 11140.846016
Rwpos46_36 in46 sp36 11140.846016
Rwpos46_37 in46 sp37 3183.098862
Rwpos46_38 in46 sp38 11140.846016
Rwpos46_39 in46 sp39 3183.098862
Rwpos46_40 in46 sp40 3183.098862
Rwpos46_41 in46 sp41 11140.846016
Rwpos46_42 in46 sp42 11140.846016
Rwpos46_43 in46 sp43 11140.846016
Rwpos46_44 in46 sp44 11140.846016
Rwpos46_45 in46 sp45 11140.846016
Rwpos46_46 in46 sp46 11140.846016
Rwpos46_47 in46 sp47 3183.098862
Rwpos46_48 in46 sp48 11140.846016
Rwpos46_49 in46 sp49 11140.846016
Rwpos46_50 in46 sp50 11140.846016
Rwpos46_51 in46 sp51 11140.846016
Rwpos46_52 in46 sp52 11140.846016
Rwpos46_53 in46 sp53 3183.098862
Rwpos46_54 in46 sp54 3183.098862
Rwpos46_55 in46 sp55 3183.098862
Rwpos46_56 in46 sp56 11140.846016
Rwpos46_57 in46 sp57 11140.846016
Rwpos46_58 in46 sp58 11140.846016
Rwpos46_59 in46 sp59 3183.098862
Rwpos46_60 in46 sp60 3183.098862
Rwpos46_61 in46 sp61 11140.846016
Rwpos46_62 in46 sp62 11140.846016
Rwpos46_63 in46 sp63 3183.098862
Rwpos46_64 in46 sp64 11140.846016
Rwpos46_65 in46 sp65 11140.846016
Rwpos46_66 in46 sp66 11140.846016
Rwpos46_67 in46 sp67 3183.098862
Rwpos46_68 in46 sp68 11140.846016
Rwpos46_69 in46 sp69 3183.098862
Rwpos46_70 in46 sp70 11140.846016
Rwpos46_71 in46 sp71 11140.846016
Rwpos46_72 in46 sp72 11140.846016
Rwpos46_73 in46 sp73 3183.098862
Rwpos46_74 in46 sp74 11140.846016
Rwpos46_75 in46 sp75 11140.846016
Rwpos46_76 in46 sp76 11140.846016
Rwpos46_77 in46 sp77 3183.098862
Rwpos46_78 in46 sp78 11140.846016
Rwpos46_79 in46 sp79 11140.846016
Rwpos46_80 in46 sp80 11140.846016
Rwpos46_81 in46 sp81 3183.098862
Rwpos46_82 in46 sp82 3183.098862
Rwpos46_83 in46 sp83 3183.098862
Rwpos46_84 in46 sp84 11140.846016
Rwpos46_85 in46 sp85 11140.846016
Rwpos46_86 in46 sp86 11140.846016
Rwpos46_87 in46 sp87 3183.098862
Rwpos46_88 in46 sp88 3183.098862
Rwpos46_89 in46 sp89 11140.846016
Rwpos46_90 in46 sp90 3183.098862
Rwpos46_91 in46 sp91 11140.846016
Rwpos46_92 in46 sp92 3183.098862
Rwpos46_93 in46 sp93 11140.846016
Rwpos46_94 in46 sp94 3183.098862
Rwpos46_95 in46 sp95 3183.098862
Rwpos46_96 in46 sp96 3183.098862
Rwpos46_97 in46 sp97 3183.098862
Rwpos46_98 in46 sp98 3183.098862
Rwpos46_99 in46 sp99 3183.098862
Rwpos46_100 in46 sp100 3183.098862
Rwpos47_1 in47 sp1 3183.098862
Rwpos47_2 in47 sp2 11140.846016
Rwpos47_3 in47 sp3 3183.098862
Rwpos47_4 in47 sp4 3183.098862
Rwpos47_5 in47 sp5 11140.846016
Rwpos47_6 in47 sp6 11140.846016
Rwpos47_7 in47 sp7 3183.098862
Rwpos47_8 in47 sp8 11140.846016
Rwpos47_9 in47 sp9 3183.098862
Rwpos47_10 in47 sp10 11140.846016
Rwpos47_11 in47 sp11 3183.098862
Rwpos47_12 in47 sp12 11140.846016
Rwpos47_13 in47 sp13 3183.098862
Rwpos47_14 in47 sp14 3183.098862
Rwpos47_15 in47 sp15 11140.846016
Rwpos47_16 in47 sp16 11140.846016
Rwpos47_17 in47 sp17 11140.846016
Rwpos47_18 in47 sp18 3183.098862
Rwpos47_19 in47 sp19 3183.098862
Rwpos47_20 in47 sp20 3183.098862
Rwpos47_21 in47 sp21 11140.846016
Rwpos47_22 in47 sp22 11140.846016
Rwpos47_23 in47 sp23 3183.098862
Rwpos47_24 in47 sp24 3183.098862
Rwpos47_25 in47 sp25 3183.098862
Rwpos47_26 in47 sp26 3183.098862
Rwpos47_27 in47 sp27 11140.846016
Rwpos47_28 in47 sp28 11140.846016
Rwpos47_29 in47 sp29 11140.846016
Rwpos47_30 in47 sp30 3183.098862
Rwpos47_31 in47 sp31 3183.098862
Rwpos47_32 in47 sp32 3183.098862
Rwpos47_33 in47 sp33 11140.846016
Rwpos47_34 in47 sp34 3183.098862
Rwpos47_35 in47 sp35 3183.098862
Rwpos47_36 in47 sp36 11140.846016
Rwpos47_37 in47 sp37 11140.846016
Rwpos47_38 in47 sp38 11140.846016
Rwpos47_39 in47 sp39 11140.846016
Rwpos47_40 in47 sp40 3183.098862
Rwpos47_41 in47 sp41 3183.098862
Rwpos47_42 in47 sp42 11140.846016
Rwpos47_43 in47 sp43 3183.098862
Rwpos47_44 in47 sp44 11140.846016
Rwpos47_45 in47 sp45 3183.098862
Rwpos47_46 in47 sp46 3183.098862
Rwpos47_47 in47 sp47 3183.098862
Rwpos47_48 in47 sp48 11140.846016
Rwpos47_49 in47 sp49 11140.846016
Rwpos47_50 in47 sp50 3183.098862
Rwpos47_51 in47 sp51 3183.098862
Rwpos47_52 in47 sp52 3183.098862
Rwpos47_53 in47 sp53 11140.846016
Rwpos47_54 in47 sp54 3183.098862
Rwpos47_55 in47 sp55 3183.098862
Rwpos47_56 in47 sp56 3183.098862
Rwpos47_57 in47 sp57 3183.098862
Rwpos47_58 in47 sp58 3183.098862
Rwpos47_59 in47 sp59 11140.846016
Rwpos47_60 in47 sp60 3183.098862
Rwpos47_61 in47 sp61 11140.846016
Rwpos47_62 in47 sp62 3183.098862
Rwpos47_63 in47 sp63 11140.846016
Rwpos47_64 in47 sp64 3183.098862
Rwpos47_65 in47 sp65 11140.846016
Rwpos47_66 in47 sp66 3183.098862
Rwpos47_67 in47 sp67 3183.098862
Rwpos47_68 in47 sp68 3183.098862
Rwpos47_69 in47 sp69 11140.846016
Rwpos47_70 in47 sp70 3183.098862
Rwpos47_71 in47 sp71 11140.846016
Rwpos47_72 in47 sp72 3183.098862
Rwpos47_73 in47 sp73 3183.098862
Rwpos47_74 in47 sp74 3183.098862
Rwpos47_75 in47 sp75 3183.098862
Rwpos47_76 in47 sp76 11140.846016
Rwpos47_77 in47 sp77 11140.846016
Rwpos47_78 in47 sp78 3183.098862
Rwpos47_79 in47 sp79 3183.098862
Rwpos47_80 in47 sp80 11140.846016
Rwpos47_81 in47 sp81 11140.846016
Rwpos47_82 in47 sp82 3183.098862
Rwpos47_83 in47 sp83 3183.098862
Rwpos47_84 in47 sp84 3183.098862
Rwpos47_85 in47 sp85 11140.846016
Rwpos47_86 in47 sp86 3183.098862
Rwpos47_87 in47 sp87 11140.846016
Rwpos47_88 in47 sp88 3183.098862
Rwpos47_89 in47 sp89 11140.846016
Rwpos47_90 in47 sp90 3183.098862
Rwpos47_91 in47 sp91 3183.098862
Rwpos47_92 in47 sp92 11140.846016
Rwpos47_93 in47 sp93 3183.098862
Rwpos47_94 in47 sp94 11140.846016
Rwpos47_95 in47 sp95 3183.098862
Rwpos47_96 in47 sp96 3183.098862
Rwpos47_97 in47 sp97 11140.846016
Rwpos47_98 in47 sp98 3183.098862
Rwpos47_99 in47 sp99 3183.098862
Rwpos47_100 in47 sp100 3183.098862
Rwpos48_1 in48 sp1 11140.846016
Rwpos48_2 in48 sp2 3183.098862
Rwpos48_3 in48 sp3 11140.846016
Rwpos48_4 in48 sp4 3183.098862
Rwpos48_5 in48 sp5 11140.846016
Rwpos48_6 in48 sp6 3183.098862
Rwpos48_7 in48 sp7 11140.846016
Rwpos48_8 in48 sp8 11140.846016
Rwpos48_9 in48 sp9 3183.098862
Rwpos48_10 in48 sp10 3183.098862
Rwpos48_11 in48 sp11 11140.846016
Rwpos48_12 in48 sp12 3183.098862
Rwpos48_13 in48 sp13 11140.846016
Rwpos48_14 in48 sp14 3183.098862
Rwpos48_15 in48 sp15 3183.098862
Rwpos48_16 in48 sp16 3183.098862
Rwpos48_17 in48 sp17 3183.098862
Rwpos48_18 in48 sp18 11140.846016
Rwpos48_19 in48 sp19 11140.846016
Rwpos48_20 in48 sp20 3183.098862
Rwpos48_21 in48 sp21 11140.846016
Rwpos48_22 in48 sp22 3183.098862
Rwpos48_23 in48 sp23 3183.098862
Rwpos48_24 in48 sp24 11140.846016
Rwpos48_25 in48 sp25 3183.098862
Rwpos48_26 in48 sp26 3183.098862
Rwpos48_27 in48 sp27 11140.846016
Rwpos48_28 in48 sp28 11140.846016
Rwpos48_29 in48 sp29 3183.098862
Rwpos48_30 in48 sp30 3183.098862
Rwpos48_31 in48 sp31 11140.846016
Rwpos48_32 in48 sp32 3183.098862
Rwpos48_33 in48 sp33 3183.098862
Rwpos48_34 in48 sp34 3183.098862
Rwpos48_35 in48 sp35 11140.846016
Rwpos48_36 in48 sp36 3183.098862
Rwpos48_37 in48 sp37 11140.846016
Rwpos48_38 in48 sp38 3183.098862
Rwpos48_39 in48 sp39 3183.098862
Rwpos48_40 in48 sp40 11140.846016
Rwpos48_41 in48 sp41 11140.846016
Rwpos48_42 in48 sp42 3183.098862
Rwpos48_43 in48 sp43 11140.846016
Rwpos48_44 in48 sp44 3183.098862
Rwpos48_45 in48 sp45 3183.098862
Rwpos48_46 in48 sp46 3183.098862
Rwpos48_47 in48 sp47 11140.846016
Rwpos48_48 in48 sp48 3183.098862
Rwpos48_49 in48 sp49 3183.098862
Rwpos48_50 in48 sp50 11140.846016
Rwpos48_51 in48 sp51 11140.846016
Rwpos48_52 in48 sp52 3183.098862
Rwpos48_53 in48 sp53 11140.846016
Rwpos48_54 in48 sp54 11140.846016
Rwpos48_55 in48 sp55 3183.098862
Rwpos48_56 in48 sp56 11140.846016
Rwpos48_57 in48 sp57 11140.846016
Rwpos48_58 in48 sp58 3183.098862
Rwpos48_59 in48 sp59 3183.098862
Rwpos48_60 in48 sp60 11140.846016
Rwpos48_61 in48 sp61 3183.098862
Rwpos48_62 in48 sp62 3183.098862
Rwpos48_63 in48 sp63 11140.846016
Rwpos48_64 in48 sp64 11140.846016
Rwpos48_65 in48 sp65 3183.098862
Rwpos48_66 in48 sp66 3183.098862
Rwpos48_67 in48 sp67 11140.846016
Rwpos48_68 in48 sp68 3183.098862
Rwpos48_69 in48 sp69 11140.846016
Rwpos48_70 in48 sp70 11140.846016
Rwpos48_71 in48 sp71 3183.098862
Rwpos48_72 in48 sp72 11140.846016
Rwpos48_73 in48 sp73 3183.098862
Rwpos48_74 in48 sp74 3183.098862
Rwpos48_75 in48 sp75 3183.098862
Rwpos48_76 in48 sp76 3183.098862
Rwpos48_77 in48 sp77 3183.098862
Rwpos48_78 in48 sp78 11140.846016
Rwpos48_79 in48 sp79 11140.846016
Rwpos48_80 in48 sp80 11140.846016
Rwpos48_81 in48 sp81 3183.098862
Rwpos48_82 in48 sp82 11140.846016
Rwpos48_83 in48 sp83 11140.846016
Rwpos48_84 in48 sp84 3183.098862
Rwpos48_85 in48 sp85 11140.846016
Rwpos48_86 in48 sp86 3183.098862
Rwpos48_87 in48 sp87 3183.098862
Rwpos48_88 in48 sp88 11140.846016
Rwpos48_89 in48 sp89 11140.846016
Rwpos48_90 in48 sp90 3183.098862
Rwpos48_91 in48 sp91 3183.098862
Rwpos48_92 in48 sp92 11140.846016
Rwpos48_93 in48 sp93 3183.098862
Rwpos48_94 in48 sp94 3183.098862
Rwpos48_95 in48 sp95 3183.098862
Rwpos48_96 in48 sp96 11140.846016
Rwpos48_97 in48 sp97 3183.098862
Rwpos48_98 in48 sp98 11140.846016
Rwpos48_99 in48 sp99 11140.846016
Rwpos48_100 in48 sp100 3183.098862
Rwpos49_1 in49 sp1 11140.846016
Rwpos49_2 in49 sp2 11140.846016
Rwpos49_3 in49 sp3 11140.846016
Rwpos49_4 in49 sp4 3183.098862
Rwpos49_5 in49 sp5 11140.846016
Rwpos49_6 in49 sp6 3183.098862
Rwpos49_7 in49 sp7 3183.098862
Rwpos49_8 in49 sp8 11140.846016
Rwpos49_9 in49 sp9 3183.098862
Rwpos49_10 in49 sp10 3183.098862
Rwpos49_11 in49 sp11 11140.846016
Rwpos49_12 in49 sp12 11140.846016
Rwpos49_13 in49 sp13 3183.098862
Rwpos49_14 in49 sp14 3183.098862
Rwpos49_15 in49 sp15 11140.846016
Rwpos49_16 in49 sp16 3183.098862
Rwpos49_17 in49 sp17 11140.846016
Rwpos49_18 in49 sp18 11140.846016
Rwpos49_19 in49 sp19 11140.846016
Rwpos49_20 in49 sp20 11140.846016
Rwpos49_21 in49 sp21 3183.098862
Rwpos49_22 in49 sp22 3183.098862
Rwpos49_23 in49 sp23 3183.098862
Rwpos49_24 in49 sp24 3183.098862
Rwpos49_25 in49 sp25 3183.098862
Rwpos49_26 in49 sp26 3183.098862
Rwpos49_27 in49 sp27 3183.098862
Rwpos49_28 in49 sp28 11140.846016
Rwpos49_29 in49 sp29 3183.098862
Rwpos49_30 in49 sp30 11140.846016
Rwpos49_31 in49 sp31 11140.846016
Rwpos49_32 in49 sp32 11140.846016
Rwpos49_33 in49 sp33 11140.846016
Rwpos49_34 in49 sp34 11140.846016
Rwpos49_35 in49 sp35 3183.098862
Rwpos49_36 in49 sp36 11140.846016
Rwpos49_37 in49 sp37 3183.098862
Rwpos49_38 in49 sp38 3183.098862
Rwpos49_39 in49 sp39 3183.098862
Rwpos49_40 in49 sp40 3183.098862
Rwpos49_41 in49 sp41 3183.098862
Rwpos49_42 in49 sp42 3183.098862
Rwpos49_43 in49 sp43 3183.098862
Rwpos49_44 in49 sp44 11140.846016
Rwpos49_45 in49 sp45 11140.846016
Rwpos49_46 in49 sp46 11140.846016
Rwpos49_47 in49 sp47 11140.846016
Rwpos49_48 in49 sp48 3183.098862
Rwpos49_49 in49 sp49 3183.098862
Rwpos49_50 in49 sp50 11140.846016
Rwpos49_51 in49 sp51 3183.098862
Rwpos49_52 in49 sp52 11140.846016
Rwpos49_53 in49 sp53 3183.098862
Rwpos49_54 in49 sp54 3183.098862
Rwpos49_55 in49 sp55 3183.098862
Rwpos49_56 in49 sp56 3183.098862
Rwpos49_57 in49 sp57 11140.846016
Rwpos49_58 in49 sp58 11140.846016
Rwpos49_59 in49 sp59 3183.098862
Rwpos49_60 in49 sp60 11140.846016
Rwpos49_61 in49 sp61 11140.846016
Rwpos49_62 in49 sp62 11140.846016
Rwpos49_63 in49 sp63 11140.846016
Rwpos49_64 in49 sp64 3183.098862
Rwpos49_65 in49 sp65 11140.846016
Rwpos49_66 in49 sp66 11140.846016
Rwpos49_67 in49 sp67 3183.098862
Rwpos49_68 in49 sp68 3183.098862
Rwpos49_69 in49 sp69 3183.098862
Rwpos49_70 in49 sp70 3183.098862
Rwpos49_71 in49 sp71 11140.846016
Rwpos49_72 in49 sp72 3183.098862
Rwpos49_73 in49 sp73 11140.846016
Rwpos49_74 in49 sp74 3183.098862
Rwpos49_75 in49 sp75 11140.846016
Rwpos49_76 in49 sp76 11140.846016
Rwpos49_77 in49 sp77 11140.846016
Rwpos49_78 in49 sp78 3183.098862
Rwpos49_79 in49 sp79 11140.846016
Rwpos49_80 in49 sp80 3183.098862
Rwpos49_81 in49 sp81 11140.846016
Rwpos49_82 in49 sp82 11140.846016
Rwpos49_83 in49 sp83 11140.846016
Rwpos49_84 in49 sp84 3183.098862
Rwpos49_85 in49 sp85 11140.846016
Rwpos49_86 in49 sp86 11140.846016
Rwpos49_87 in49 sp87 3183.098862
Rwpos49_88 in49 sp88 3183.098862
Rwpos49_89 in49 sp89 11140.846016
Rwpos49_90 in49 sp90 3183.098862
Rwpos49_91 in49 sp91 3183.098862
Rwpos49_92 in49 sp92 3183.098862
Rwpos49_93 in49 sp93 11140.846016
Rwpos49_94 in49 sp94 3183.098862
Rwpos49_95 in49 sp95 3183.098862
Rwpos49_96 in49 sp96 3183.098862
Rwpos49_97 in49 sp97 3183.098862
Rwpos49_98 in49 sp98 11140.846016
Rwpos49_99 in49 sp99 3183.098862
Rwpos49_100 in49 sp100 11140.846016
Rwpos50_1 in50 sp1 3183.098862
Rwpos50_2 in50 sp2 11140.846016
Rwpos50_3 in50 sp3 3183.098862
Rwpos50_4 in50 sp4 3183.098862
Rwpos50_5 in50 sp5 11140.846016
Rwpos50_6 in50 sp6 3183.098862
Rwpos50_7 in50 sp7 11140.846016
Rwpos50_8 in50 sp8 11140.846016
Rwpos50_9 in50 sp9 11140.846016
Rwpos50_10 in50 sp10 3183.098862
Rwpos50_11 in50 sp11 11140.846016
Rwpos50_12 in50 sp12 3183.098862
Rwpos50_13 in50 sp13 11140.846016
Rwpos50_14 in50 sp14 11140.846016
Rwpos50_15 in50 sp15 11140.846016
Rwpos50_16 in50 sp16 3183.098862
Rwpos50_17 in50 sp17 3183.098862
Rwpos50_18 in50 sp18 3183.098862
Rwpos50_19 in50 sp19 3183.098862
Rwpos50_20 in50 sp20 11140.846016
Rwpos50_21 in50 sp21 11140.846016
Rwpos50_22 in50 sp22 11140.846016
Rwpos50_23 in50 sp23 3183.098862
Rwpos50_24 in50 sp24 11140.846016
Rwpos50_25 in50 sp25 3183.098862
Rwpos50_26 in50 sp26 3183.098862
Rwpos50_27 in50 sp27 11140.846016
Rwpos50_28 in50 sp28 3183.098862
Rwpos50_29 in50 sp29 3183.098862
Rwpos50_30 in50 sp30 11140.846016
Rwpos50_31 in50 sp31 11140.846016
Rwpos50_32 in50 sp32 11140.846016
Rwpos50_33 in50 sp33 3183.098862
Rwpos50_34 in50 sp34 11140.846016
Rwpos50_35 in50 sp35 11140.846016
Rwpos50_36 in50 sp36 3183.098862
Rwpos50_37 in50 sp37 11140.846016
Rwpos50_38 in50 sp38 11140.846016
Rwpos50_39 in50 sp39 3183.098862
Rwpos50_40 in50 sp40 3183.098862
Rwpos50_41 in50 sp41 3183.098862
Rwpos50_42 in50 sp42 3183.098862
Rwpos50_43 in50 sp43 11140.846016
Rwpos50_44 in50 sp44 11140.846016
Rwpos50_45 in50 sp45 3183.098862
Rwpos50_46 in50 sp46 11140.846016
Rwpos50_47 in50 sp47 3183.098862
Rwpos50_48 in50 sp48 11140.846016
Rwpos50_49 in50 sp49 11140.846016
Rwpos50_50 in50 sp50 3183.098862
Rwpos50_51 in50 sp51 11140.846016
Rwpos50_52 in50 sp52 3183.098862
Rwpos50_53 in50 sp53 3183.098862
Rwpos50_54 in50 sp54 3183.098862
Rwpos50_55 in50 sp55 11140.846016
Rwpos50_56 in50 sp56 3183.098862
Rwpos50_57 in50 sp57 3183.098862
Rwpos50_58 in50 sp58 3183.098862
Rwpos50_59 in50 sp59 3183.098862
Rwpos50_60 in50 sp60 11140.846016
Rwpos50_61 in50 sp61 3183.098862
Rwpos50_62 in50 sp62 11140.846016
Rwpos50_63 in50 sp63 11140.846016
Rwpos50_64 in50 sp64 3183.098862
Rwpos50_65 in50 sp65 3183.098862
Rwpos50_66 in50 sp66 11140.846016
Rwpos50_67 in50 sp67 3183.098862
Rwpos50_68 in50 sp68 11140.846016
Rwpos50_69 in50 sp69 3183.098862
Rwpos50_70 in50 sp70 3183.098862
Rwpos50_71 in50 sp71 3183.098862
Rwpos50_72 in50 sp72 3183.098862
Rwpos50_73 in50 sp73 11140.846016
Rwpos50_74 in50 sp74 3183.098862
Rwpos50_75 in50 sp75 11140.846016
Rwpos50_76 in50 sp76 3183.098862
Rwpos50_77 in50 sp77 11140.846016
Rwpos50_78 in50 sp78 11140.846016
Rwpos50_79 in50 sp79 3183.098862
Rwpos50_80 in50 sp80 11140.846016
Rwpos50_81 in50 sp81 3183.098862
Rwpos50_82 in50 sp82 11140.846016
Rwpos50_83 in50 sp83 3183.098862
Rwpos50_84 in50 sp84 11140.846016
Rwpos50_85 in50 sp85 11140.846016
Rwpos50_86 in50 sp86 3183.098862
Rwpos50_87 in50 sp87 11140.846016
Rwpos50_88 in50 sp88 11140.846016
Rwpos50_89 in50 sp89 3183.098862
Rwpos50_90 in50 sp90 11140.846016
Rwpos50_91 in50 sp91 11140.846016
Rwpos50_92 in50 sp92 11140.846016
Rwpos50_93 in50 sp93 11140.846016
Rwpos50_94 in50 sp94 11140.846016
Rwpos50_95 in50 sp95 11140.846016
Rwpos50_96 in50 sp96 11140.846016
Rwpos50_97 in50 sp97 3183.098862
Rwpos50_98 in50 sp98 3183.098862
Rwpos50_99 in50 sp99 11140.846016
Rwpos50_100 in50 sp100 3183.098862
Rwpos51_1 in51 sp1 11140.846016
Rwpos51_2 in51 sp2 11140.846016
Rwpos51_3 in51 sp3 11140.846016
Rwpos51_4 in51 sp4 3183.098862
Rwpos51_5 in51 sp5 3183.098862
Rwpos51_6 in51 sp6 11140.846016
Rwpos51_7 in51 sp7 3183.098862
Rwpos51_8 in51 sp8 3183.098862
Rwpos51_9 in51 sp9 3183.098862
Rwpos51_10 in51 sp10 11140.846016
Rwpos51_11 in51 sp11 11140.846016
Rwpos51_12 in51 sp12 3183.098862
Rwpos51_13 in51 sp13 11140.846016
Rwpos51_14 in51 sp14 3183.098862
Rwpos51_15 in51 sp15 3183.098862
Rwpos51_16 in51 sp16 3183.098862
Rwpos51_17 in51 sp17 3183.098862
Rwpos51_18 in51 sp18 3183.098862
Rwpos51_19 in51 sp19 3183.098862
Rwpos51_20 in51 sp20 3183.098862
Rwpos51_21 in51 sp21 11140.846016
Rwpos51_22 in51 sp22 11140.846016
Rwpos51_23 in51 sp23 11140.846016
Rwpos51_24 in51 sp24 3183.098862
Rwpos51_25 in51 sp25 3183.098862
Rwpos51_26 in51 sp26 11140.846016
Rwpos51_27 in51 sp27 11140.846016
Rwpos51_28 in51 sp28 11140.846016
Rwpos51_29 in51 sp29 11140.846016
Rwpos51_30 in51 sp30 3183.098862
Rwpos51_31 in51 sp31 11140.846016
Rwpos51_32 in51 sp32 11140.846016
Rwpos51_33 in51 sp33 11140.846016
Rwpos51_34 in51 sp34 3183.098862
Rwpos51_35 in51 sp35 3183.098862
Rwpos51_36 in51 sp36 3183.098862
Rwpos51_37 in51 sp37 3183.098862
Rwpos51_38 in51 sp38 11140.846016
Rwpos51_39 in51 sp39 11140.846016
Rwpos51_40 in51 sp40 3183.098862
Rwpos51_41 in51 sp41 3183.098862
Rwpos51_42 in51 sp42 3183.098862
Rwpos51_43 in51 sp43 11140.846016
Rwpos51_44 in51 sp44 11140.846016
Rwpos51_45 in51 sp45 11140.846016
Rwpos51_46 in51 sp46 3183.098862
Rwpos51_47 in51 sp47 3183.098862
Rwpos51_48 in51 sp48 11140.846016
Rwpos51_49 in51 sp49 11140.846016
Rwpos51_50 in51 sp50 11140.846016
Rwpos51_51 in51 sp51 3183.098862
Rwpos51_52 in51 sp52 3183.098862
Rwpos51_53 in51 sp53 11140.846016
Rwpos51_54 in51 sp54 11140.846016
Rwpos51_55 in51 sp55 11140.846016
Rwpos51_56 in51 sp56 3183.098862
Rwpos51_57 in51 sp57 3183.098862
Rwpos51_58 in51 sp58 3183.098862
Rwpos51_59 in51 sp59 11140.846016
Rwpos51_60 in51 sp60 3183.098862
Rwpos51_61 in51 sp61 3183.098862
Rwpos51_62 in51 sp62 3183.098862
Rwpos51_63 in51 sp63 3183.098862
Rwpos51_64 in51 sp64 11140.846016
Rwpos51_65 in51 sp65 11140.846016
Rwpos51_66 in51 sp66 11140.846016
Rwpos51_67 in51 sp67 3183.098862
Rwpos51_68 in51 sp68 3183.098862
Rwpos51_69 in51 sp69 11140.846016
Rwpos51_70 in51 sp70 11140.846016
Rwpos51_71 in51 sp71 3183.098862
Rwpos51_72 in51 sp72 3183.098862
Rwpos51_73 in51 sp73 3183.098862
Rwpos51_74 in51 sp74 3183.098862
Rwpos51_75 in51 sp75 11140.846016
Rwpos51_76 in51 sp76 11140.846016
Rwpos51_77 in51 sp77 11140.846016
Rwpos51_78 in51 sp78 3183.098862
Rwpos51_79 in51 sp79 11140.846016
Rwpos51_80 in51 sp80 11140.846016
Rwpos51_81 in51 sp81 3183.098862
Rwpos51_82 in51 sp82 11140.846016
Rwpos51_83 in51 sp83 3183.098862
Rwpos51_84 in51 sp84 3183.098862
Rwpos51_85 in51 sp85 11140.846016
Rwpos51_86 in51 sp86 11140.846016
Rwpos51_87 in51 sp87 3183.098862
Rwpos51_88 in51 sp88 3183.098862
Rwpos51_89 in51 sp89 3183.098862
Rwpos51_90 in51 sp90 11140.846016
Rwpos51_91 in51 sp91 11140.846016
Rwpos51_92 in51 sp92 3183.098862
Rwpos51_93 in51 sp93 11140.846016
Rwpos51_94 in51 sp94 3183.098862
Rwpos51_95 in51 sp95 3183.098862
Rwpos51_96 in51 sp96 3183.098862
Rwpos51_97 in51 sp97 11140.846016
Rwpos51_98 in51 sp98 11140.846016
Rwpos51_99 in51 sp99 3183.098862
Rwpos51_100 in51 sp100 3183.098862
Rwpos52_1 in52 sp1 11140.846016
Rwpos52_2 in52 sp2 11140.846016
Rwpos52_3 in52 sp3 11140.846016
Rwpos52_4 in52 sp4 3183.098862
Rwpos52_5 in52 sp5 3183.098862
Rwpos52_6 in52 sp6 11140.846016
Rwpos52_7 in52 sp7 3183.098862
Rwpos52_8 in52 sp8 3183.098862
Rwpos52_9 in52 sp9 11140.846016
Rwpos52_10 in52 sp10 3183.098862
Rwpos52_11 in52 sp11 11140.846016
Rwpos52_12 in52 sp12 11140.846016
Rwpos52_13 in52 sp13 11140.846016
Rwpos52_14 in52 sp14 11140.846016
Rwpos52_15 in52 sp15 3183.098862
Rwpos52_16 in52 sp16 3183.098862
Rwpos52_17 in52 sp17 11140.846016
Rwpos52_18 in52 sp18 3183.098862
Rwpos52_19 in52 sp19 3183.098862
Rwpos52_20 in52 sp20 3183.098862
Rwpos52_21 in52 sp21 3183.098862
Rwpos52_22 in52 sp22 11140.846016
Rwpos52_23 in52 sp23 11140.846016
Rwpos52_24 in52 sp24 3183.098862
Rwpos52_25 in52 sp25 3183.098862
Rwpos52_26 in52 sp26 3183.098862
Rwpos52_27 in52 sp27 3183.098862
Rwpos52_28 in52 sp28 11140.846016
Rwpos52_29 in52 sp29 11140.846016
Rwpos52_30 in52 sp30 11140.846016
Rwpos52_31 in52 sp31 3183.098862
Rwpos52_32 in52 sp32 3183.098862
Rwpos52_33 in52 sp33 11140.846016
Rwpos52_34 in52 sp34 11140.846016
Rwpos52_35 in52 sp35 11140.846016
Rwpos52_36 in52 sp36 3183.098862
Rwpos52_37 in52 sp37 11140.846016
Rwpos52_38 in52 sp38 11140.846016
Rwpos52_39 in52 sp39 3183.098862
Rwpos52_40 in52 sp40 11140.846016
Rwpos52_41 in52 sp41 11140.846016
Rwpos52_42 in52 sp42 11140.846016
Rwpos52_43 in52 sp43 11140.846016
Rwpos52_44 in52 sp44 3183.098862
Rwpos52_45 in52 sp45 11140.846016
Rwpos52_46 in52 sp46 3183.098862
Rwpos52_47 in52 sp47 3183.098862
Rwpos52_48 in52 sp48 3183.098862
Rwpos52_49 in52 sp49 11140.846016
Rwpos52_50 in52 sp50 3183.098862
Rwpos52_51 in52 sp51 3183.098862
Rwpos52_52 in52 sp52 3183.098862
Rwpos52_53 in52 sp53 11140.846016
Rwpos52_54 in52 sp54 3183.098862
Rwpos52_55 in52 sp55 3183.098862
Rwpos52_56 in52 sp56 11140.846016
Rwpos52_57 in52 sp57 11140.846016
Rwpos52_58 in52 sp58 11140.846016
Rwpos52_59 in52 sp59 11140.846016
Rwpos52_60 in52 sp60 3183.098862
Rwpos52_61 in52 sp61 3183.098862
Rwpos52_62 in52 sp62 3183.098862
Rwpos52_63 in52 sp63 3183.098862
Rwpos52_64 in52 sp64 3183.098862
Rwpos52_65 in52 sp65 3183.098862
Rwpos52_66 in52 sp66 11140.846016
Rwpos52_67 in52 sp67 3183.098862
Rwpos52_68 in52 sp68 3183.098862
Rwpos52_69 in52 sp69 11140.846016
Rwpos52_70 in52 sp70 3183.098862
Rwpos52_71 in52 sp71 11140.846016
Rwpos52_72 in52 sp72 11140.846016
Rwpos52_73 in52 sp73 11140.846016
Rwpos52_74 in52 sp74 11140.846016
Rwpos52_75 in52 sp75 11140.846016
Rwpos52_76 in52 sp76 11140.846016
Rwpos52_77 in52 sp77 3183.098862
Rwpos52_78 in52 sp78 3183.098862
Rwpos52_79 in52 sp79 11140.846016
Rwpos52_80 in52 sp80 3183.098862
Rwpos52_81 in52 sp81 3183.098862
Rwpos52_82 in52 sp82 11140.846016
Rwpos52_83 in52 sp83 3183.098862
Rwpos52_84 in52 sp84 3183.098862
Rwpos52_85 in52 sp85 11140.846016
Rwpos52_86 in52 sp86 11140.846016
Rwpos52_87 in52 sp87 3183.098862
Rwpos52_88 in52 sp88 11140.846016
Rwpos52_89 in52 sp89 11140.846016
Rwpos52_90 in52 sp90 11140.846016
Rwpos52_91 in52 sp91 3183.098862
Rwpos52_92 in52 sp92 11140.846016
Rwpos52_93 in52 sp93 3183.098862
Rwpos52_94 in52 sp94 11140.846016
Rwpos52_95 in52 sp95 11140.846016
Rwpos52_96 in52 sp96 3183.098862
Rwpos52_97 in52 sp97 3183.098862
Rwpos52_98 in52 sp98 3183.098862
Rwpos52_99 in52 sp99 11140.846016
Rwpos52_100 in52 sp100 3183.098862
Rwpos53_1 in53 sp1 11140.846016
Rwpos53_2 in53 sp2 11140.846016
Rwpos53_3 in53 sp3 11140.846016
Rwpos53_4 in53 sp4 3183.098862
Rwpos53_5 in53 sp5 3183.098862
Rwpos53_6 in53 sp6 3183.098862
Rwpos53_7 in53 sp7 3183.098862
Rwpos53_8 in53 sp8 11140.846016
Rwpos53_9 in53 sp9 3183.098862
Rwpos53_10 in53 sp10 3183.098862
Rwpos53_11 in53 sp11 11140.846016
Rwpos53_12 in53 sp12 3183.098862
Rwpos53_13 in53 sp13 3183.098862
Rwpos53_14 in53 sp14 3183.098862
Rwpos53_15 in53 sp15 11140.846016
Rwpos53_16 in53 sp16 3183.098862
Rwpos53_17 in53 sp17 11140.846016
Rwpos53_18 in53 sp18 11140.846016
Rwpos53_19 in53 sp19 11140.846016
Rwpos53_20 in53 sp20 11140.846016
Rwpos53_21 in53 sp21 11140.846016
Rwpos53_22 in53 sp22 11140.846016
Rwpos53_23 in53 sp23 3183.098862
Rwpos53_24 in53 sp24 11140.846016
Rwpos53_25 in53 sp25 3183.098862
Rwpos53_26 in53 sp26 11140.846016
Rwpos53_27 in53 sp27 3183.098862
Rwpos53_28 in53 sp28 11140.846016
Rwpos53_29 in53 sp29 3183.098862
Rwpos53_30 in53 sp30 3183.098862
Rwpos53_31 in53 sp31 11140.846016
Rwpos53_32 in53 sp32 11140.846016
Rwpos53_33 in53 sp33 11140.846016
Rwpos53_34 in53 sp34 11140.846016
Rwpos53_35 in53 sp35 11140.846016
Rwpos53_36 in53 sp36 3183.098862
Rwpos53_37 in53 sp37 3183.098862
Rwpos53_38 in53 sp38 3183.098862
Rwpos53_39 in53 sp39 3183.098862
Rwpos53_40 in53 sp40 11140.846016
Rwpos53_41 in53 sp41 3183.098862
Rwpos53_42 in53 sp42 3183.098862
Rwpos53_43 in53 sp43 11140.846016
Rwpos53_44 in53 sp44 11140.846016
Rwpos53_45 in53 sp45 3183.098862
Rwpos53_46 in53 sp46 11140.846016
Rwpos53_47 in53 sp47 11140.846016
Rwpos53_48 in53 sp48 3183.098862
Rwpos53_49 in53 sp49 11140.846016
Rwpos53_50 in53 sp50 3183.098862
Rwpos53_51 in53 sp51 11140.846016
Rwpos53_52 in53 sp52 11140.846016
Rwpos53_53 in53 sp53 11140.846016
Rwpos53_54 in53 sp54 3183.098862
Rwpos53_55 in53 sp55 3183.098862
Rwpos53_56 in53 sp56 11140.846016
Rwpos53_57 in53 sp57 3183.098862
Rwpos53_58 in53 sp58 3183.098862
Rwpos53_59 in53 sp59 11140.846016
Rwpos53_60 in53 sp60 11140.846016
Rwpos53_61 in53 sp61 3183.098862
Rwpos53_62 in53 sp62 11140.846016
Rwpos53_63 in53 sp63 11140.846016
Rwpos53_64 in53 sp64 3183.098862
Rwpos53_65 in53 sp65 3183.098862
Rwpos53_66 in53 sp66 11140.846016
Rwpos53_67 in53 sp67 11140.846016
Rwpos53_68 in53 sp68 3183.098862
Rwpos53_69 in53 sp69 3183.098862
Rwpos53_70 in53 sp70 3183.098862
Rwpos53_71 in53 sp71 3183.098862
Rwpos53_72 in53 sp72 11140.846016
Rwpos53_73 in53 sp73 3183.098862
Rwpos53_74 in53 sp74 3183.098862
Rwpos53_75 in53 sp75 3183.098862
Rwpos53_76 in53 sp76 11140.846016
Rwpos53_77 in53 sp77 3183.098862
Rwpos53_78 in53 sp78 11140.846016
Rwpos53_79 in53 sp79 11140.846016
Rwpos53_80 in53 sp80 3183.098862
Rwpos53_81 in53 sp81 3183.098862
Rwpos53_82 in53 sp82 11140.846016
Rwpos53_83 in53 sp83 11140.846016
Rwpos53_84 in53 sp84 11140.846016
Rwpos53_85 in53 sp85 11140.846016
Rwpos53_86 in53 sp86 3183.098862
Rwpos53_87 in53 sp87 3183.098862
Rwpos53_88 in53 sp88 11140.846016
Rwpos53_89 in53 sp89 3183.098862
Rwpos53_90 in53 sp90 11140.846016
Rwpos53_91 in53 sp91 3183.098862
Rwpos53_92 in53 sp92 3183.098862
Rwpos53_93 in53 sp93 3183.098862
Rwpos53_94 in53 sp94 11140.846016
Rwpos53_95 in53 sp95 11140.846016
Rwpos53_96 in53 sp96 3183.098862
Rwpos53_97 in53 sp97 3183.098862
Rwpos53_98 in53 sp98 11140.846016
Rwpos53_99 in53 sp99 3183.098862
Rwpos53_100 in53 sp100 3183.098862
Rwpos54_1 in54 sp1 3183.098862
Rwpos54_2 in54 sp2 11140.846016
Rwpos54_3 in54 sp3 11140.846016
Rwpos54_4 in54 sp4 3183.098862
Rwpos54_5 in54 sp5 3183.098862
Rwpos54_6 in54 sp6 3183.098862
Rwpos54_7 in54 sp7 3183.098862
Rwpos54_8 in54 sp8 11140.846016
Rwpos54_9 in54 sp9 11140.846016
Rwpos54_10 in54 sp10 11140.846016
Rwpos54_11 in54 sp11 11140.846016
Rwpos54_12 in54 sp12 3183.098862
Rwpos54_13 in54 sp13 11140.846016
Rwpos54_14 in54 sp14 11140.846016
Rwpos54_15 in54 sp15 11140.846016
Rwpos54_16 in54 sp16 11140.846016
Rwpos54_17 in54 sp17 11140.846016
Rwpos54_18 in54 sp18 11140.846016
Rwpos54_19 in54 sp19 11140.846016
Rwpos54_20 in54 sp20 3183.098862
Rwpos54_21 in54 sp21 3183.098862
Rwpos54_22 in54 sp22 3183.098862
Rwpos54_23 in54 sp23 11140.846016
Rwpos54_24 in54 sp24 11140.846016
Rwpos54_25 in54 sp25 3183.098862
Rwpos54_26 in54 sp26 3183.098862
Rwpos54_27 in54 sp27 11140.846016
Rwpos54_28 in54 sp28 11140.846016
Rwpos54_29 in54 sp29 3183.098862
Rwpos54_30 in54 sp30 3183.098862
Rwpos54_31 in54 sp31 3183.098862
Rwpos54_32 in54 sp32 11140.846016
Rwpos54_33 in54 sp33 3183.098862
Rwpos54_34 in54 sp34 3183.098862
Rwpos54_35 in54 sp35 3183.098862
Rwpos54_36 in54 sp36 3183.098862
Rwpos54_37 in54 sp37 11140.846016
Rwpos54_38 in54 sp38 11140.846016
Rwpos54_39 in54 sp39 11140.846016
Rwpos54_40 in54 sp40 3183.098862
Rwpos54_41 in54 sp41 11140.846016
Rwpos54_42 in54 sp42 11140.846016
Rwpos54_43 in54 sp43 3183.098862
Rwpos54_44 in54 sp44 11140.846016
Rwpos54_45 in54 sp45 11140.846016
Rwpos54_46 in54 sp46 3183.098862
Rwpos54_47 in54 sp47 3183.098862
Rwpos54_48 in54 sp48 3183.098862
Rwpos54_49 in54 sp49 3183.098862
Rwpos54_50 in54 sp50 11140.846016
Rwpos54_51 in54 sp51 3183.098862
Rwpos54_52 in54 sp52 3183.098862
Rwpos54_53 in54 sp53 11140.846016
Rwpos54_54 in54 sp54 3183.098862
Rwpos54_55 in54 sp55 11140.846016
Rwpos54_56 in54 sp56 11140.846016
Rwpos54_57 in54 sp57 3183.098862
Rwpos54_58 in54 sp58 11140.846016
Rwpos54_59 in54 sp59 3183.098862
Rwpos54_60 in54 sp60 3183.098862
Rwpos54_61 in54 sp61 11140.846016
Rwpos54_62 in54 sp62 3183.098862
Rwpos54_63 in54 sp63 11140.846016
Rwpos54_64 in54 sp64 11140.846016
Rwpos54_65 in54 sp65 11140.846016
Rwpos54_66 in54 sp66 11140.846016
Rwpos54_67 in54 sp67 11140.846016
Rwpos54_68 in54 sp68 3183.098862
Rwpos54_69 in54 sp69 11140.846016
Rwpos54_70 in54 sp70 11140.846016
Rwpos54_71 in54 sp71 3183.098862
Rwpos54_72 in54 sp72 3183.098862
Rwpos54_73 in54 sp73 3183.098862
Rwpos54_74 in54 sp74 3183.098862
Rwpos54_75 in54 sp75 11140.846016
Rwpos54_76 in54 sp76 11140.846016
Rwpos54_77 in54 sp77 11140.846016
Rwpos54_78 in54 sp78 11140.846016
Rwpos54_79 in54 sp79 3183.098862
Rwpos54_80 in54 sp80 11140.846016
Rwpos54_81 in54 sp81 11140.846016
Rwpos54_82 in54 sp82 3183.098862
Rwpos54_83 in54 sp83 11140.846016
Rwpos54_84 in54 sp84 3183.098862
Rwpos54_85 in54 sp85 3183.098862
Rwpos54_86 in54 sp86 3183.098862
Rwpos54_87 in54 sp87 11140.846016
Rwpos54_88 in54 sp88 11140.846016
Rwpos54_89 in54 sp89 11140.846016
Rwpos54_90 in54 sp90 11140.846016
Rwpos54_91 in54 sp91 3183.098862
Rwpos54_92 in54 sp92 3183.098862
Rwpos54_93 in54 sp93 11140.846016
Rwpos54_94 in54 sp94 3183.098862
Rwpos54_95 in54 sp95 11140.846016
Rwpos54_96 in54 sp96 11140.846016
Rwpos54_97 in54 sp97 3183.098862
Rwpos54_98 in54 sp98 3183.098862
Rwpos54_99 in54 sp99 11140.846016
Rwpos54_100 in54 sp100 11140.846016
Rwpos55_1 in55 sp1 11140.846016
Rwpos55_2 in55 sp2 3183.098862
Rwpos55_3 in55 sp3 11140.846016
Rwpos55_4 in55 sp4 11140.846016
Rwpos55_5 in55 sp5 3183.098862
Rwpos55_6 in55 sp6 11140.846016
Rwpos55_7 in55 sp7 11140.846016
Rwpos55_8 in55 sp8 3183.098862
Rwpos55_9 in55 sp9 3183.098862
Rwpos55_10 in55 sp10 11140.846016
Rwpos55_11 in55 sp11 11140.846016
Rwpos55_12 in55 sp12 11140.846016
Rwpos55_13 in55 sp13 3183.098862
Rwpos55_14 in55 sp14 3183.098862
Rwpos55_15 in55 sp15 11140.846016
Rwpos55_16 in55 sp16 11140.846016
Rwpos55_17 in55 sp17 11140.846016
Rwpos55_18 in55 sp18 11140.846016
Rwpos55_19 in55 sp19 11140.846016
Rwpos55_20 in55 sp20 3183.098862
Rwpos55_21 in55 sp21 11140.846016
Rwpos55_22 in55 sp22 3183.098862
Rwpos55_23 in55 sp23 11140.846016
Rwpos55_24 in55 sp24 3183.098862
Rwpos55_25 in55 sp25 11140.846016
Rwpos55_26 in55 sp26 11140.846016
Rwpos55_27 in55 sp27 3183.098862
Rwpos55_28 in55 sp28 3183.098862
Rwpos55_29 in55 sp29 3183.098862
Rwpos55_30 in55 sp30 11140.846016
Rwpos55_31 in55 sp31 3183.098862
Rwpos55_32 in55 sp32 11140.846016
Rwpos55_33 in55 sp33 11140.846016
Rwpos55_34 in55 sp34 11140.846016
Rwpos55_35 in55 sp35 3183.098862
Rwpos55_36 in55 sp36 11140.846016
Rwpos55_37 in55 sp37 11140.846016
Rwpos55_38 in55 sp38 3183.098862
Rwpos55_39 in55 sp39 3183.098862
Rwpos55_40 in55 sp40 11140.846016
Rwpos55_41 in55 sp41 11140.846016
Rwpos55_42 in55 sp42 11140.846016
Rwpos55_43 in55 sp43 3183.098862
Rwpos55_44 in55 sp44 11140.846016
Rwpos55_45 in55 sp45 11140.846016
Rwpos55_46 in55 sp46 11140.846016
Rwpos55_47 in55 sp47 3183.098862
Rwpos55_48 in55 sp48 11140.846016
Rwpos55_49 in55 sp49 3183.098862
Rwpos55_50 in55 sp50 3183.098862
Rwpos55_51 in55 sp51 11140.846016
Rwpos55_52 in55 sp52 11140.846016
Rwpos55_53 in55 sp53 11140.846016
Rwpos55_54 in55 sp54 3183.098862
Rwpos55_55 in55 sp55 3183.098862
Rwpos55_56 in55 sp56 11140.846016
Rwpos55_57 in55 sp57 11140.846016
Rwpos55_58 in55 sp58 3183.098862
Rwpos55_59 in55 sp59 11140.846016
Rwpos55_60 in55 sp60 11140.846016
Rwpos55_61 in55 sp61 11140.846016
Rwpos55_62 in55 sp62 11140.846016
Rwpos55_63 in55 sp63 11140.846016
Rwpos55_64 in55 sp64 11140.846016
Rwpos55_65 in55 sp65 3183.098862
Rwpos55_66 in55 sp66 11140.846016
Rwpos55_67 in55 sp67 3183.098862
Rwpos55_68 in55 sp68 3183.098862
Rwpos55_69 in55 sp69 11140.846016
Rwpos55_70 in55 sp70 3183.098862
Rwpos55_71 in55 sp71 11140.846016
Rwpos55_72 in55 sp72 3183.098862
Rwpos55_73 in55 sp73 3183.098862
Rwpos55_74 in55 sp74 11140.846016
Rwpos55_75 in55 sp75 11140.846016
Rwpos55_76 in55 sp76 11140.846016
Rwpos55_77 in55 sp77 3183.098862
Rwpos55_78 in55 sp78 11140.846016
Rwpos55_79 in55 sp79 11140.846016
Rwpos55_80 in55 sp80 11140.846016
Rwpos55_81 in55 sp81 11140.846016
Rwpos55_82 in55 sp82 11140.846016
Rwpos55_83 in55 sp83 3183.098862
Rwpos55_84 in55 sp84 3183.098862
Rwpos55_85 in55 sp85 11140.846016
Rwpos55_86 in55 sp86 11140.846016
Rwpos55_87 in55 sp87 3183.098862
Rwpos55_88 in55 sp88 3183.098862
Rwpos55_89 in55 sp89 3183.098862
Rwpos55_90 in55 sp90 3183.098862
Rwpos55_91 in55 sp91 11140.846016
Rwpos55_92 in55 sp92 3183.098862
Rwpos55_93 in55 sp93 11140.846016
Rwpos55_94 in55 sp94 3183.098862
Rwpos55_95 in55 sp95 3183.098862
Rwpos55_96 in55 sp96 11140.846016
Rwpos55_97 in55 sp97 11140.846016
Rwpos55_98 in55 sp98 3183.098862
Rwpos55_99 in55 sp99 3183.098862
Rwpos55_100 in55 sp100 3183.098862
Rwpos56_1 in56 sp1 11140.846016
Rwpos56_2 in56 sp2 3183.098862
Rwpos56_3 in56 sp3 3183.098862
Rwpos56_4 in56 sp4 3183.098862
Rwpos56_5 in56 sp5 3183.098862
Rwpos56_6 in56 sp6 11140.846016
Rwpos56_7 in56 sp7 11140.846016
Rwpos56_8 in56 sp8 3183.098862
Rwpos56_9 in56 sp9 11140.846016
Rwpos56_10 in56 sp10 11140.846016
Rwpos56_11 in56 sp11 11140.846016
Rwpos56_12 in56 sp12 11140.846016
Rwpos56_13 in56 sp13 11140.846016
Rwpos56_14 in56 sp14 11140.846016
Rwpos56_15 in56 sp15 3183.098862
Rwpos56_16 in56 sp16 3183.098862
Rwpos56_17 in56 sp17 11140.846016
Rwpos56_18 in56 sp18 3183.098862
Rwpos56_19 in56 sp19 11140.846016
Rwpos56_20 in56 sp20 3183.098862
Rwpos56_21 in56 sp21 3183.098862
Rwpos56_22 in56 sp22 3183.098862
Rwpos56_23 in56 sp23 11140.846016
Rwpos56_24 in56 sp24 3183.098862
Rwpos56_25 in56 sp25 3183.098862
Rwpos56_26 in56 sp26 3183.098862
Rwpos56_27 in56 sp27 11140.846016
Rwpos56_28 in56 sp28 11140.846016
Rwpos56_29 in56 sp29 11140.846016
Rwpos56_30 in56 sp30 11140.846016
Rwpos56_31 in56 sp31 3183.098862
Rwpos56_32 in56 sp32 3183.098862
Rwpos56_33 in56 sp33 11140.846016
Rwpos56_34 in56 sp34 3183.098862
Rwpos56_35 in56 sp35 11140.846016
Rwpos56_36 in56 sp36 3183.098862
Rwpos56_37 in56 sp37 3183.098862
Rwpos56_38 in56 sp38 3183.098862
Rwpos56_39 in56 sp39 3183.098862
Rwpos56_40 in56 sp40 3183.098862
Rwpos56_41 in56 sp41 3183.098862
Rwpos56_42 in56 sp42 11140.846016
Rwpos56_43 in56 sp43 3183.098862
Rwpos56_44 in56 sp44 11140.846016
Rwpos56_45 in56 sp45 11140.846016
Rwpos56_46 in56 sp46 11140.846016
Rwpos56_47 in56 sp47 3183.098862
Rwpos56_48 in56 sp48 3183.098862
Rwpos56_49 in56 sp49 11140.846016
Rwpos56_50 in56 sp50 11140.846016
Rwpos56_51 in56 sp51 3183.098862
Rwpos56_52 in56 sp52 3183.098862
Rwpos56_53 in56 sp53 3183.098862
Rwpos56_54 in56 sp54 11140.846016
Rwpos56_55 in56 sp55 11140.846016
Rwpos56_56 in56 sp56 3183.098862
Rwpos56_57 in56 sp57 11140.846016
Rwpos56_58 in56 sp58 11140.846016
Rwpos56_59 in56 sp59 3183.098862
Rwpos56_60 in56 sp60 11140.846016
Rwpos56_61 in56 sp61 11140.846016
Rwpos56_62 in56 sp62 11140.846016
Rwpos56_63 in56 sp63 3183.098862
Rwpos56_64 in56 sp64 3183.098862
Rwpos56_65 in56 sp65 11140.846016
Rwpos56_66 in56 sp66 3183.098862
Rwpos56_67 in56 sp67 3183.098862
Rwpos56_68 in56 sp68 3183.098862
Rwpos56_69 in56 sp69 3183.098862
Rwpos56_70 in56 sp70 11140.846016
Rwpos56_71 in56 sp71 3183.098862
Rwpos56_72 in56 sp72 3183.098862
Rwpos56_73 in56 sp73 3183.098862
Rwpos56_74 in56 sp74 11140.846016
Rwpos56_75 in56 sp75 3183.098862
Rwpos56_76 in56 sp76 11140.846016
Rwpos56_77 in56 sp77 11140.846016
Rwpos56_78 in56 sp78 11140.846016
Rwpos56_79 in56 sp79 3183.098862
Rwpos56_80 in56 sp80 3183.098862
Rwpos56_81 in56 sp81 11140.846016
Rwpos56_82 in56 sp82 3183.098862
Rwpos56_83 in56 sp83 3183.098862
Rwpos56_84 in56 sp84 3183.098862
Rwpos56_85 in56 sp85 11140.846016
Rwpos56_86 in56 sp86 11140.846016
Rwpos56_87 in56 sp87 11140.846016
Rwpos56_88 in56 sp88 3183.098862
Rwpos56_89 in56 sp89 3183.098862
Rwpos56_90 in56 sp90 11140.846016
Rwpos56_91 in56 sp91 11140.846016
Rwpos56_92 in56 sp92 3183.098862
Rwpos56_93 in56 sp93 11140.846016
Rwpos56_94 in56 sp94 11140.846016
Rwpos56_95 in56 sp95 3183.098862
Rwpos56_96 in56 sp96 3183.098862
Rwpos56_97 in56 sp97 11140.846016
Rwpos56_98 in56 sp98 11140.846016
Rwpos56_99 in56 sp99 3183.098862
Rwpos56_100 in56 sp100 3183.098862
Rwpos57_1 in57 sp1 3183.098862
Rwpos57_2 in57 sp2 11140.846016
Rwpos57_3 in57 sp3 11140.846016
Rwpos57_4 in57 sp4 11140.846016
Rwpos57_5 in57 sp5 3183.098862
Rwpos57_6 in57 sp6 11140.846016
Rwpos57_7 in57 sp7 11140.846016
Rwpos57_8 in57 sp8 3183.098862
Rwpos57_9 in57 sp9 3183.098862
Rwpos57_10 in57 sp10 3183.098862
Rwpos57_11 in57 sp11 3183.098862
Rwpos57_12 in57 sp12 3183.098862
Rwpos57_13 in57 sp13 11140.846016
Rwpos57_14 in57 sp14 11140.846016
Rwpos57_15 in57 sp15 3183.098862
Rwpos57_16 in57 sp16 3183.098862
Rwpos57_17 in57 sp17 11140.846016
Rwpos57_18 in57 sp18 11140.846016
Rwpos57_19 in57 sp19 11140.846016
Rwpos57_20 in57 sp20 11140.846016
Rwpos57_21 in57 sp21 3183.098862
Rwpos57_22 in57 sp22 11140.846016
Rwpos57_23 in57 sp23 11140.846016
Rwpos57_24 in57 sp24 11140.846016
Rwpos57_25 in57 sp25 3183.098862
Rwpos57_26 in57 sp26 3183.098862
Rwpos57_27 in57 sp27 3183.098862
Rwpos57_28 in57 sp28 3183.098862
Rwpos57_29 in57 sp29 3183.098862
Rwpos57_30 in57 sp30 11140.846016
Rwpos57_31 in57 sp31 3183.098862
Rwpos57_32 in57 sp32 3183.098862
Rwpos57_33 in57 sp33 11140.846016
Rwpos57_34 in57 sp34 11140.846016
Rwpos57_35 in57 sp35 11140.846016
Rwpos57_36 in57 sp36 3183.098862
Rwpos57_37 in57 sp37 3183.098862
Rwpos57_38 in57 sp38 11140.846016
Rwpos57_39 in57 sp39 3183.098862
Rwpos57_40 in57 sp40 11140.846016
Rwpos57_41 in57 sp41 3183.098862
Rwpos57_42 in57 sp42 11140.846016
Rwpos57_43 in57 sp43 11140.846016
Rwpos57_44 in57 sp44 3183.098862
Rwpos57_45 in57 sp45 3183.098862
Rwpos57_46 in57 sp46 11140.846016
Rwpos57_47 in57 sp47 3183.098862
Rwpos57_48 in57 sp48 3183.098862
Rwpos57_49 in57 sp49 11140.846016
Rwpos57_50 in57 sp50 11140.846016
Rwpos57_51 in57 sp51 3183.098862
Rwpos57_52 in57 sp52 11140.846016
Rwpos57_53 in57 sp53 11140.846016
Rwpos57_54 in57 sp54 11140.846016
Rwpos57_55 in57 sp55 3183.098862
Rwpos57_56 in57 sp56 11140.846016
Rwpos57_57 in57 sp57 3183.098862
Rwpos57_58 in57 sp58 3183.098862
Rwpos57_59 in57 sp59 11140.846016
Rwpos57_60 in57 sp60 3183.098862
Rwpos57_61 in57 sp61 3183.098862
Rwpos57_62 in57 sp62 3183.098862
Rwpos57_63 in57 sp63 11140.846016
Rwpos57_64 in57 sp64 3183.098862
Rwpos57_65 in57 sp65 3183.098862
Rwpos57_66 in57 sp66 3183.098862
Rwpos57_67 in57 sp67 11140.846016
Rwpos57_68 in57 sp68 11140.846016
Rwpos57_69 in57 sp69 11140.846016
Rwpos57_70 in57 sp70 11140.846016
Rwpos57_71 in57 sp71 3183.098862
Rwpos57_72 in57 sp72 11140.846016
Rwpos57_73 in57 sp73 3183.098862
Rwpos57_74 in57 sp74 3183.098862
Rwpos57_75 in57 sp75 3183.098862
Rwpos57_76 in57 sp76 3183.098862
Rwpos57_77 in57 sp77 11140.846016
Rwpos57_78 in57 sp78 11140.846016
Rwpos57_79 in57 sp79 3183.098862
Rwpos57_80 in57 sp80 3183.098862
Rwpos57_81 in57 sp81 3183.098862
Rwpos57_82 in57 sp82 3183.098862
Rwpos57_83 in57 sp83 11140.846016
Rwpos57_84 in57 sp84 3183.098862
Rwpos57_85 in57 sp85 3183.098862
Rwpos57_86 in57 sp86 3183.098862
Rwpos57_87 in57 sp87 3183.098862
Rwpos57_88 in57 sp88 3183.098862
Rwpos57_89 in57 sp89 3183.098862
Rwpos57_90 in57 sp90 11140.846016
Rwpos57_91 in57 sp91 11140.846016
Rwpos57_92 in57 sp92 11140.846016
Rwpos57_93 in57 sp93 11140.846016
Rwpos57_94 in57 sp94 11140.846016
Rwpos57_95 in57 sp95 3183.098862
Rwpos57_96 in57 sp96 11140.846016
Rwpos57_97 in57 sp97 3183.098862
Rwpos57_98 in57 sp98 3183.098862
Rwpos57_99 in57 sp99 11140.846016
Rwpos57_100 in57 sp100 11140.846016
Rwpos58_1 in58 sp1 3183.098862
Rwpos58_2 in58 sp2 11140.846016
Rwpos58_3 in58 sp3 3183.098862
Rwpos58_4 in58 sp4 3183.098862
Rwpos58_5 in58 sp5 3183.098862
Rwpos58_6 in58 sp6 3183.098862
Rwpos58_7 in58 sp7 3183.098862
Rwpos58_8 in58 sp8 3183.098862
Rwpos58_9 in58 sp9 3183.098862
Rwpos58_10 in58 sp10 11140.846016
Rwpos58_11 in58 sp11 11140.846016
Rwpos58_12 in58 sp12 11140.846016
Rwpos58_13 in58 sp13 3183.098862
Rwpos58_14 in58 sp14 3183.098862
Rwpos58_15 in58 sp15 11140.846016
Rwpos58_16 in58 sp16 11140.846016
Rwpos58_17 in58 sp17 11140.846016
Rwpos58_18 in58 sp18 3183.098862
Rwpos58_19 in58 sp19 3183.098862
Rwpos58_20 in58 sp20 11140.846016
Rwpos58_21 in58 sp21 3183.098862
Rwpos58_22 in58 sp22 3183.098862
Rwpos58_23 in58 sp23 3183.098862
Rwpos58_24 in58 sp24 3183.098862
Rwpos58_25 in58 sp25 3183.098862
Rwpos58_26 in58 sp26 11140.846016
Rwpos58_27 in58 sp27 11140.846016
Rwpos58_28 in58 sp28 11140.846016
Rwpos58_29 in58 sp29 3183.098862
Rwpos58_30 in58 sp30 3183.098862
Rwpos58_31 in58 sp31 11140.846016
Rwpos58_32 in58 sp32 11140.846016
Rwpos58_33 in58 sp33 3183.098862
Rwpos58_34 in58 sp34 11140.846016
Rwpos58_35 in58 sp35 3183.098862
Rwpos58_36 in58 sp36 3183.098862
Rwpos58_37 in58 sp37 3183.098862
Rwpos58_38 in58 sp38 11140.846016
Rwpos58_39 in58 sp39 3183.098862
Rwpos58_40 in58 sp40 11140.846016
Rwpos58_41 in58 sp41 3183.098862
Rwpos58_42 in58 sp42 11140.846016
Rwpos58_43 in58 sp43 11140.846016
Rwpos58_44 in58 sp44 3183.098862
Rwpos58_45 in58 sp45 3183.098862
Rwpos58_46 in58 sp46 3183.098862
Rwpos58_47 in58 sp47 11140.846016
Rwpos58_48 in58 sp48 3183.098862
Rwpos58_49 in58 sp49 3183.098862
Rwpos58_50 in58 sp50 11140.846016
Rwpos58_51 in58 sp51 3183.098862
Rwpos58_52 in58 sp52 3183.098862
Rwpos58_53 in58 sp53 11140.846016
Rwpos58_54 in58 sp54 11140.846016
Rwpos58_55 in58 sp55 3183.098862
Rwpos58_56 in58 sp56 11140.846016
Rwpos58_57 in58 sp57 3183.098862
Rwpos58_58 in58 sp58 3183.098862
Rwpos58_59 in58 sp59 11140.846016
Rwpos58_60 in58 sp60 3183.098862
Rwpos58_61 in58 sp61 11140.846016
Rwpos58_62 in58 sp62 11140.846016
Rwpos58_63 in58 sp63 11140.846016
Rwpos58_64 in58 sp64 11140.846016
Rwpos58_65 in58 sp65 3183.098862
Rwpos58_66 in58 sp66 3183.098862
Rwpos58_67 in58 sp67 3183.098862
Rwpos58_68 in58 sp68 11140.846016
Rwpos58_69 in58 sp69 11140.846016
Rwpos58_70 in58 sp70 11140.846016
Rwpos58_71 in58 sp71 11140.846016
Rwpos58_72 in58 sp72 11140.846016
Rwpos58_73 in58 sp73 3183.098862
Rwpos58_74 in58 sp74 3183.098862
Rwpos58_75 in58 sp75 11140.846016
Rwpos58_76 in58 sp76 3183.098862
Rwpos58_77 in58 sp77 3183.098862
Rwpos58_78 in58 sp78 3183.098862
Rwpos58_79 in58 sp79 3183.098862
Rwpos58_80 in58 sp80 3183.098862
Rwpos58_81 in58 sp81 11140.846016
Rwpos58_82 in58 sp82 11140.846016
Rwpos58_83 in58 sp83 3183.098862
Rwpos58_84 in58 sp84 3183.098862
Rwpos58_85 in58 sp85 11140.846016
Rwpos58_86 in58 sp86 11140.846016
Rwpos58_87 in58 sp87 3183.098862
Rwpos58_88 in58 sp88 3183.098862
Rwpos58_89 in58 sp89 3183.098862
Rwpos58_90 in58 sp90 11140.846016
Rwpos58_91 in58 sp91 3183.098862
Rwpos58_92 in58 sp92 3183.098862
Rwpos58_93 in58 sp93 3183.098862
Rwpos58_94 in58 sp94 3183.098862
Rwpos58_95 in58 sp95 3183.098862
Rwpos58_96 in58 sp96 11140.846016
Rwpos58_97 in58 sp97 3183.098862
Rwpos58_98 in58 sp98 11140.846016
Rwpos58_99 in58 sp99 3183.098862
Rwpos58_100 in58 sp100 3183.098862
Rwpos59_1 in59 sp1 3183.098862
Rwpos59_2 in59 sp2 3183.098862
Rwpos59_3 in59 sp3 3183.098862
Rwpos59_4 in59 sp4 11140.846016
Rwpos59_5 in59 sp5 3183.098862
Rwpos59_6 in59 sp6 3183.098862
Rwpos59_7 in59 sp7 11140.846016
Rwpos59_8 in59 sp8 3183.098862
Rwpos59_9 in59 sp9 11140.846016
Rwpos59_10 in59 sp10 3183.098862
Rwpos59_11 in59 sp11 3183.098862
Rwpos59_12 in59 sp12 3183.098862
Rwpos59_13 in59 sp13 11140.846016
Rwpos59_14 in59 sp14 3183.098862
Rwpos59_15 in59 sp15 11140.846016
Rwpos59_16 in59 sp16 3183.098862
Rwpos59_17 in59 sp17 11140.846016
Rwpos59_18 in59 sp18 3183.098862
Rwpos59_19 in59 sp19 11140.846016
Rwpos59_20 in59 sp20 3183.098862
Rwpos59_21 in59 sp21 11140.846016
Rwpos59_22 in59 sp22 11140.846016
Rwpos59_23 in59 sp23 3183.098862
Rwpos59_24 in59 sp24 3183.098862
Rwpos59_25 in59 sp25 3183.098862
Rwpos59_26 in59 sp26 11140.846016
Rwpos59_27 in59 sp27 11140.846016
Rwpos59_28 in59 sp28 3183.098862
Rwpos59_29 in59 sp29 11140.846016
Rwpos59_30 in59 sp30 3183.098862
Rwpos59_31 in59 sp31 3183.098862
Rwpos59_32 in59 sp32 3183.098862
Rwpos59_33 in59 sp33 3183.098862
Rwpos59_34 in59 sp34 3183.098862
Rwpos59_35 in59 sp35 11140.846016
Rwpos59_36 in59 sp36 3183.098862
Rwpos59_37 in59 sp37 3183.098862
Rwpos59_38 in59 sp38 3183.098862
Rwpos59_39 in59 sp39 3183.098862
Rwpos59_40 in59 sp40 3183.098862
Rwpos59_41 in59 sp41 3183.098862
Rwpos59_42 in59 sp42 11140.846016
Rwpos59_43 in59 sp43 11140.846016
Rwpos59_44 in59 sp44 3183.098862
Rwpos59_45 in59 sp45 11140.846016
Rwpos59_46 in59 sp46 11140.846016
Rwpos59_47 in59 sp47 11140.846016
Rwpos59_48 in59 sp48 3183.098862
Rwpos59_49 in59 sp49 3183.098862
Rwpos59_50 in59 sp50 3183.098862
Rwpos59_51 in59 sp51 11140.846016
Rwpos59_52 in59 sp52 11140.846016
Rwpos59_53 in59 sp53 3183.098862
Rwpos59_54 in59 sp54 3183.098862
Rwpos59_55 in59 sp55 11140.846016
Rwpos59_56 in59 sp56 3183.098862
Rwpos59_57 in59 sp57 3183.098862
Rwpos59_58 in59 sp58 11140.846016
Rwpos59_59 in59 sp59 11140.846016
Rwpos59_60 in59 sp60 3183.098862
Rwpos59_61 in59 sp61 3183.098862
Rwpos59_62 in59 sp62 3183.098862
Rwpos59_63 in59 sp63 3183.098862
Rwpos59_64 in59 sp64 3183.098862
Rwpos59_65 in59 sp65 3183.098862
Rwpos59_66 in59 sp66 3183.098862
Rwpos59_67 in59 sp67 11140.846016
Rwpos59_68 in59 sp68 11140.846016
Rwpos59_69 in59 sp69 3183.098862
Rwpos59_70 in59 sp70 11140.846016
Rwpos59_71 in59 sp71 3183.098862
Rwpos59_72 in59 sp72 3183.098862
Rwpos59_73 in59 sp73 3183.098862
Rwpos59_74 in59 sp74 3183.098862
Rwpos59_75 in59 sp75 11140.846016
Rwpos59_76 in59 sp76 11140.846016
Rwpos59_77 in59 sp77 11140.846016
Rwpos59_78 in59 sp78 11140.846016
Rwpos59_79 in59 sp79 3183.098862
Rwpos59_80 in59 sp80 3183.098862
Rwpos59_81 in59 sp81 3183.098862
Rwpos59_82 in59 sp82 11140.846016
Rwpos59_83 in59 sp83 3183.098862
Rwpos59_84 in59 sp84 3183.098862
Rwpos59_85 in59 sp85 11140.846016
Rwpos59_86 in59 sp86 3183.098862
Rwpos59_87 in59 sp87 3183.098862
Rwpos59_88 in59 sp88 3183.098862
Rwpos59_89 in59 sp89 3183.098862
Rwpos59_90 in59 sp90 11140.846016
Rwpos59_91 in59 sp91 11140.846016
Rwpos59_92 in59 sp92 3183.098862
Rwpos59_93 in59 sp93 3183.098862
Rwpos59_94 in59 sp94 3183.098862
Rwpos59_95 in59 sp95 11140.846016
Rwpos59_96 in59 sp96 11140.846016
Rwpos59_97 in59 sp97 11140.846016
Rwpos59_98 in59 sp98 3183.098862
Rwpos59_99 in59 sp99 3183.098862
Rwpos59_100 in59 sp100 3183.098862
Rwpos60_1 in60 sp1 11140.846016
Rwpos60_2 in60 sp2 3183.098862
Rwpos60_3 in60 sp3 11140.846016
Rwpos60_4 in60 sp4 3183.098862
Rwpos60_5 in60 sp5 11140.846016
Rwpos60_6 in60 sp6 3183.098862
Rwpos60_7 in60 sp7 11140.846016
Rwpos60_8 in60 sp8 11140.846016
Rwpos60_9 in60 sp9 3183.098862
Rwpos60_10 in60 sp10 11140.846016
Rwpos60_11 in60 sp11 11140.846016
Rwpos60_12 in60 sp12 11140.846016
Rwpos60_13 in60 sp13 11140.846016
Rwpos60_14 in60 sp14 11140.846016
Rwpos60_15 in60 sp15 3183.098862
Rwpos60_16 in60 sp16 11140.846016
Rwpos60_17 in60 sp17 3183.098862
Rwpos60_18 in60 sp18 3183.098862
Rwpos60_19 in60 sp19 3183.098862
Rwpos60_20 in60 sp20 3183.098862
Rwpos60_21 in60 sp21 3183.098862
Rwpos60_22 in60 sp22 3183.098862
Rwpos60_23 in60 sp23 11140.846016
Rwpos60_24 in60 sp24 11140.846016
Rwpos60_25 in60 sp25 3183.098862
Rwpos60_26 in60 sp26 11140.846016
Rwpos60_27 in60 sp27 3183.098862
Rwpos60_28 in60 sp28 11140.846016
Rwpos60_29 in60 sp29 3183.098862
Rwpos60_30 in60 sp30 11140.846016
Rwpos60_31 in60 sp31 3183.098862
Rwpos60_32 in60 sp32 3183.098862
Rwpos60_33 in60 sp33 3183.098862
Rwpos60_34 in60 sp34 3183.098862
Rwpos60_35 in60 sp35 11140.846016
Rwpos60_36 in60 sp36 3183.098862
Rwpos60_37 in60 sp37 3183.098862
Rwpos60_38 in60 sp38 3183.098862
Rwpos60_39 in60 sp39 11140.846016
Rwpos60_40 in60 sp40 11140.846016
Rwpos60_41 in60 sp41 3183.098862
Rwpos60_42 in60 sp42 11140.846016
Rwpos60_43 in60 sp43 3183.098862
Rwpos60_44 in60 sp44 11140.846016
Rwpos60_45 in60 sp45 11140.846016
Rwpos60_46 in60 sp46 11140.846016
Rwpos60_47 in60 sp47 3183.098862
Rwpos60_48 in60 sp48 3183.098862
Rwpos60_49 in60 sp49 3183.098862
Rwpos60_50 in60 sp50 3183.098862
Rwpos60_51 in60 sp51 3183.098862
Rwpos60_52 in60 sp52 3183.098862
Rwpos60_53 in60 sp53 3183.098862
Rwpos60_54 in60 sp54 11140.846016
Rwpos60_55 in60 sp55 11140.846016
Rwpos60_56 in60 sp56 11140.846016
Rwpos60_57 in60 sp57 3183.098862
Rwpos60_58 in60 sp58 11140.846016
Rwpos60_59 in60 sp59 3183.098862
Rwpos60_60 in60 sp60 11140.846016
Rwpos60_61 in60 sp61 3183.098862
Rwpos60_62 in60 sp62 11140.846016
Rwpos60_63 in60 sp63 3183.098862
Rwpos60_64 in60 sp64 3183.098862
Rwpos60_65 in60 sp65 3183.098862
Rwpos60_66 in60 sp66 3183.098862
Rwpos60_67 in60 sp67 3183.098862
Rwpos60_68 in60 sp68 3183.098862
Rwpos60_69 in60 sp69 3183.098862
Rwpos60_70 in60 sp70 11140.846016
Rwpos60_71 in60 sp71 11140.846016
Rwpos60_72 in60 sp72 3183.098862
Rwpos60_73 in60 sp73 3183.098862
Rwpos60_74 in60 sp74 3183.098862
Rwpos60_75 in60 sp75 11140.846016
Rwpos60_76 in60 sp76 11140.846016
Rwpos60_77 in60 sp77 11140.846016
Rwpos60_78 in60 sp78 11140.846016
Rwpos60_79 in60 sp79 3183.098862
Rwpos60_80 in60 sp80 3183.098862
Rwpos60_81 in60 sp81 11140.846016
Rwpos60_82 in60 sp82 3183.098862
Rwpos60_83 in60 sp83 3183.098862
Rwpos60_84 in60 sp84 3183.098862
Rwpos60_85 in60 sp85 3183.098862
Rwpos60_86 in60 sp86 11140.846016
Rwpos60_87 in60 sp87 11140.846016
Rwpos60_88 in60 sp88 3183.098862
Rwpos60_89 in60 sp89 3183.098862
Rwpos60_90 in60 sp90 11140.846016
Rwpos60_91 in60 sp91 11140.846016
Rwpos60_92 in60 sp92 11140.846016
Rwpos60_93 in60 sp93 11140.846016
Rwpos60_94 in60 sp94 11140.846016
Rwpos60_95 in60 sp95 3183.098862
Rwpos60_96 in60 sp96 3183.098862
Rwpos60_97 in60 sp97 3183.098862
Rwpos60_98 in60 sp98 3183.098862
Rwpos60_99 in60 sp99 11140.846016
Rwpos60_100 in60 sp100 3183.098862
Rwpos61_1 in61 sp1 3183.098862
Rwpos61_2 in61 sp2 11140.846016
Rwpos61_3 in61 sp3 3183.098862
Rwpos61_4 in61 sp4 3183.098862
Rwpos61_5 in61 sp5 3183.098862
Rwpos61_6 in61 sp6 11140.846016
Rwpos61_7 in61 sp7 11140.846016
Rwpos61_8 in61 sp8 11140.846016
Rwpos61_9 in61 sp9 11140.846016
Rwpos61_10 in61 sp10 11140.846016
Rwpos61_11 in61 sp11 3183.098862
Rwpos61_12 in61 sp12 3183.098862
Rwpos61_13 in61 sp13 11140.846016
Rwpos61_14 in61 sp14 3183.098862
Rwpos61_15 in61 sp15 3183.098862
Rwpos61_16 in61 sp16 3183.098862
Rwpos61_17 in61 sp17 3183.098862
Rwpos61_18 in61 sp18 11140.846016
Rwpos61_19 in61 sp19 11140.846016
Rwpos61_20 in61 sp20 3183.098862
Rwpos61_21 in61 sp21 3183.098862
Rwpos61_22 in61 sp22 11140.846016
Rwpos61_23 in61 sp23 3183.098862
Rwpos61_24 in61 sp24 3183.098862
Rwpos61_25 in61 sp25 11140.846016
Rwpos61_26 in61 sp26 11140.846016
Rwpos61_27 in61 sp27 11140.846016
Rwpos61_28 in61 sp28 3183.098862
Rwpos61_29 in61 sp29 11140.846016
Rwpos61_30 in61 sp30 3183.098862
Rwpos61_31 in61 sp31 3183.098862
Rwpos61_32 in61 sp32 3183.098862
Rwpos61_33 in61 sp33 11140.846016
Rwpos61_34 in61 sp34 11140.846016
Rwpos61_35 in61 sp35 11140.846016
Rwpos61_36 in61 sp36 3183.098862
Rwpos61_37 in61 sp37 3183.098862
Rwpos61_38 in61 sp38 11140.846016
Rwpos61_39 in61 sp39 11140.846016
Rwpos61_40 in61 sp40 3183.098862
Rwpos61_41 in61 sp41 3183.098862
Rwpos61_42 in61 sp42 11140.846016
Rwpos61_43 in61 sp43 11140.846016
Rwpos61_44 in61 sp44 3183.098862
Rwpos61_45 in61 sp45 11140.846016
Rwpos61_46 in61 sp46 11140.846016
Rwpos61_47 in61 sp47 3183.098862
Rwpos61_48 in61 sp48 3183.098862
Rwpos61_49 in61 sp49 3183.098862
Rwpos61_50 in61 sp50 3183.098862
Rwpos61_51 in61 sp51 11140.846016
Rwpos61_52 in61 sp52 11140.846016
Rwpos61_53 in61 sp53 3183.098862
Rwpos61_54 in61 sp54 11140.846016
Rwpos61_55 in61 sp55 11140.846016
Rwpos61_56 in61 sp56 11140.846016
Rwpos61_57 in61 sp57 3183.098862
Rwpos61_58 in61 sp58 3183.098862
Rwpos61_59 in61 sp59 3183.098862
Rwpos61_60 in61 sp60 3183.098862
Rwpos61_61 in61 sp61 11140.846016
Rwpos61_62 in61 sp62 11140.846016
Rwpos61_63 in61 sp63 3183.098862
Rwpos61_64 in61 sp64 3183.098862
Rwpos61_65 in61 sp65 3183.098862
Rwpos61_66 in61 sp66 11140.846016
Rwpos61_67 in61 sp67 11140.846016
Rwpos61_68 in61 sp68 3183.098862
Rwpos61_69 in61 sp69 3183.098862
Rwpos61_70 in61 sp70 11140.846016
Rwpos61_71 in61 sp71 11140.846016
Rwpos61_72 in61 sp72 11140.846016
Rwpos61_73 in61 sp73 3183.098862
Rwpos61_74 in61 sp74 3183.098862
Rwpos61_75 in61 sp75 3183.098862
Rwpos61_76 in61 sp76 3183.098862
Rwpos61_77 in61 sp77 3183.098862
Rwpos61_78 in61 sp78 11140.846016
Rwpos61_79 in61 sp79 3183.098862
Rwpos61_80 in61 sp80 3183.098862
Rwpos61_81 in61 sp81 11140.846016
Rwpos61_82 in61 sp82 3183.098862
Rwpos61_83 in61 sp83 11140.846016
Rwpos61_84 in61 sp84 3183.098862
Rwpos61_85 in61 sp85 3183.098862
Rwpos61_86 in61 sp86 11140.846016
Rwpos61_87 in61 sp87 3183.098862
Rwpos61_88 in61 sp88 11140.846016
Rwpos61_89 in61 sp89 3183.098862
Rwpos61_90 in61 sp90 11140.846016
Rwpos61_91 in61 sp91 3183.098862
Rwpos61_92 in61 sp92 3183.098862
Rwpos61_93 in61 sp93 11140.846016
Rwpos61_94 in61 sp94 3183.098862
Rwpos61_95 in61 sp95 3183.098862
Rwpos61_96 in61 sp96 3183.098862
Rwpos61_97 in61 sp97 3183.098862
Rwpos61_98 in61 sp98 3183.098862
Rwpos61_99 in61 sp99 11140.846016
Rwpos61_100 in61 sp100 3183.098862
Rwpos62_1 in62 sp1 11140.846016
Rwpos62_2 in62 sp2 11140.846016
Rwpos62_3 in62 sp3 3183.098862
Rwpos62_4 in62 sp4 11140.846016
Rwpos62_5 in62 sp5 3183.098862
Rwpos62_6 in62 sp6 11140.846016
Rwpos62_7 in62 sp7 11140.846016
Rwpos62_8 in62 sp8 3183.098862
Rwpos62_9 in62 sp9 3183.098862
Rwpos62_10 in62 sp10 3183.098862
Rwpos62_11 in62 sp11 3183.098862
Rwpos62_12 in62 sp12 3183.098862
Rwpos62_13 in62 sp13 3183.098862
Rwpos62_14 in62 sp14 3183.098862
Rwpos62_15 in62 sp15 11140.846016
Rwpos62_16 in62 sp16 3183.098862
Rwpos62_17 in62 sp17 11140.846016
Rwpos62_18 in62 sp18 3183.098862
Rwpos62_19 in62 sp19 3183.098862
Rwpos62_20 in62 sp20 11140.846016
Rwpos62_21 in62 sp21 3183.098862
Rwpos62_22 in62 sp22 11140.846016
Rwpos62_23 in62 sp23 3183.098862
Rwpos62_24 in62 sp24 3183.098862
Rwpos62_25 in62 sp25 11140.846016
Rwpos62_26 in62 sp26 11140.846016
Rwpos62_27 in62 sp27 3183.098862
Rwpos62_28 in62 sp28 11140.846016
Rwpos62_29 in62 sp29 3183.098862
Rwpos62_30 in62 sp30 3183.098862
Rwpos62_31 in62 sp31 11140.846016
Rwpos62_32 in62 sp32 11140.846016
Rwpos62_33 in62 sp33 11140.846016
Rwpos62_34 in62 sp34 11140.846016
Rwpos62_35 in62 sp35 3183.098862
Rwpos62_36 in62 sp36 11140.846016
Rwpos62_37 in62 sp37 3183.098862
Rwpos62_38 in62 sp38 3183.098862
Rwpos62_39 in62 sp39 11140.846016
Rwpos62_40 in62 sp40 3183.098862
Rwpos62_41 in62 sp41 3183.098862
Rwpos62_42 in62 sp42 3183.098862
Rwpos62_43 in62 sp43 3183.098862
Rwpos62_44 in62 sp44 3183.098862
Rwpos62_45 in62 sp45 3183.098862
Rwpos62_46 in62 sp46 11140.846016
Rwpos62_47 in62 sp47 11140.846016
Rwpos62_48 in62 sp48 3183.098862
Rwpos62_49 in62 sp49 3183.098862
Rwpos62_50 in62 sp50 3183.098862
Rwpos62_51 in62 sp51 3183.098862
Rwpos62_52 in62 sp52 11140.846016
Rwpos62_53 in62 sp53 3183.098862
Rwpos62_54 in62 sp54 3183.098862
Rwpos62_55 in62 sp55 3183.098862
Rwpos62_56 in62 sp56 11140.846016
Rwpos62_57 in62 sp57 3183.098862
Rwpos62_58 in62 sp58 3183.098862
Rwpos62_59 in62 sp59 3183.098862
Rwpos62_60 in62 sp60 11140.846016
Rwpos62_61 in62 sp61 3183.098862
Rwpos62_62 in62 sp62 11140.846016
Rwpos62_63 in62 sp63 11140.846016
Rwpos62_64 in62 sp64 3183.098862
Rwpos62_65 in62 sp65 3183.098862
Rwpos62_66 in62 sp66 11140.846016
Rwpos62_67 in62 sp67 3183.098862
Rwpos62_68 in62 sp68 3183.098862
Rwpos62_69 in62 sp69 11140.846016
Rwpos62_70 in62 sp70 11140.846016
Rwpos62_71 in62 sp71 3183.098862
Rwpos62_72 in62 sp72 11140.846016
Rwpos62_73 in62 sp73 3183.098862
Rwpos62_74 in62 sp74 3183.098862
Rwpos62_75 in62 sp75 11140.846016
Rwpos62_76 in62 sp76 3183.098862
Rwpos62_77 in62 sp77 3183.098862
Rwpos62_78 in62 sp78 11140.846016
Rwpos62_79 in62 sp79 3183.098862
Rwpos62_80 in62 sp80 11140.846016
Rwpos62_81 in62 sp81 11140.846016
Rwpos62_82 in62 sp82 11140.846016
Rwpos62_83 in62 sp83 3183.098862
Rwpos62_84 in62 sp84 3183.098862
Rwpos62_85 in62 sp85 11140.846016
Rwpos62_86 in62 sp86 11140.846016
Rwpos62_87 in62 sp87 3183.098862
Rwpos62_88 in62 sp88 3183.098862
Rwpos62_89 in62 sp89 3183.098862
Rwpos62_90 in62 sp90 3183.098862
Rwpos62_91 in62 sp91 11140.846016
Rwpos62_92 in62 sp92 11140.846016
Rwpos62_93 in62 sp93 3183.098862
Rwpos62_94 in62 sp94 3183.098862
Rwpos62_95 in62 sp95 11140.846016
Rwpos62_96 in62 sp96 3183.098862
Rwpos62_97 in62 sp97 11140.846016
Rwpos62_98 in62 sp98 11140.846016
Rwpos62_99 in62 sp99 3183.098862
Rwpos62_100 in62 sp100 3183.098862
Rwpos63_1 in63 sp1 3183.098862
Rwpos63_2 in63 sp2 11140.846016
Rwpos63_3 in63 sp3 3183.098862
Rwpos63_4 in63 sp4 11140.846016
Rwpos63_5 in63 sp5 3183.098862
Rwpos63_6 in63 sp6 3183.098862
Rwpos63_7 in63 sp7 11140.846016
Rwpos63_8 in63 sp8 11140.846016
Rwpos63_9 in63 sp9 11140.846016
Rwpos63_10 in63 sp10 3183.098862
Rwpos63_11 in63 sp11 11140.846016
Rwpos63_12 in63 sp12 3183.098862
Rwpos63_13 in63 sp13 3183.098862
Rwpos63_14 in63 sp14 3183.098862
Rwpos63_15 in63 sp15 3183.098862
Rwpos63_16 in63 sp16 3183.098862
Rwpos63_17 in63 sp17 11140.846016
Rwpos63_18 in63 sp18 11140.846016
Rwpos63_19 in63 sp19 3183.098862
Rwpos63_20 in63 sp20 11140.846016
Rwpos63_21 in63 sp21 3183.098862
Rwpos63_22 in63 sp22 3183.098862
Rwpos63_23 in63 sp23 3183.098862
Rwpos63_24 in63 sp24 11140.846016
Rwpos63_25 in63 sp25 3183.098862
Rwpos63_26 in63 sp26 11140.846016
Rwpos63_27 in63 sp27 11140.846016
Rwpos63_28 in63 sp28 3183.098862
Rwpos63_29 in63 sp29 3183.098862
Rwpos63_30 in63 sp30 3183.098862
Rwpos63_31 in63 sp31 11140.846016
Rwpos63_32 in63 sp32 11140.846016
Rwpos63_33 in63 sp33 11140.846016
Rwpos63_34 in63 sp34 3183.098862
Rwpos63_35 in63 sp35 3183.098862
Rwpos63_36 in63 sp36 3183.098862
Rwpos63_37 in63 sp37 11140.846016
Rwpos63_38 in63 sp38 3183.098862
Rwpos63_39 in63 sp39 11140.846016
Rwpos63_40 in63 sp40 3183.098862
Rwpos63_41 in63 sp41 11140.846016
Rwpos63_42 in63 sp42 11140.846016
Rwpos63_43 in63 sp43 11140.846016
Rwpos63_44 in63 sp44 3183.098862
Rwpos63_45 in63 sp45 11140.846016
Rwpos63_46 in63 sp46 11140.846016
Rwpos63_47 in63 sp47 11140.846016
Rwpos63_48 in63 sp48 3183.098862
Rwpos63_49 in63 sp49 3183.098862
Rwpos63_50 in63 sp50 3183.098862
Rwpos63_51 in63 sp51 3183.098862
Rwpos63_52 in63 sp52 11140.846016
Rwpos63_53 in63 sp53 3183.098862
Rwpos63_54 in63 sp54 3183.098862
Rwpos63_55 in63 sp55 11140.846016
Rwpos63_56 in63 sp56 11140.846016
Rwpos63_57 in63 sp57 3183.098862
Rwpos63_58 in63 sp58 3183.098862
Rwpos63_59 in63 sp59 3183.098862
Rwpos63_60 in63 sp60 11140.846016
Rwpos63_61 in63 sp61 11140.846016
Rwpos63_62 in63 sp62 3183.098862
Rwpos63_63 in63 sp63 11140.846016
Rwpos63_64 in63 sp64 11140.846016
Rwpos63_65 in63 sp65 11140.846016
Rwpos63_66 in63 sp66 11140.846016
Rwpos63_67 in63 sp67 11140.846016
Rwpos63_68 in63 sp68 3183.098862
Rwpos63_69 in63 sp69 11140.846016
Rwpos63_70 in63 sp70 11140.846016
Rwpos63_71 in63 sp71 3183.098862
Rwpos63_72 in63 sp72 3183.098862
Rwpos63_73 in63 sp73 3183.098862
Rwpos63_74 in63 sp74 3183.098862
Rwpos63_75 in63 sp75 3183.098862
Rwpos63_76 in63 sp76 3183.098862
Rwpos63_77 in63 sp77 3183.098862
Rwpos63_78 in63 sp78 11140.846016
Rwpos63_79 in63 sp79 3183.098862
Rwpos63_80 in63 sp80 3183.098862
Rwpos63_81 in63 sp81 11140.846016
Rwpos63_82 in63 sp82 3183.098862
Rwpos63_83 in63 sp83 3183.098862
Rwpos63_84 in63 sp84 3183.098862
Rwpos63_85 in63 sp85 3183.098862
Rwpos63_86 in63 sp86 11140.846016
Rwpos63_87 in63 sp87 3183.098862
Rwpos63_88 in63 sp88 3183.098862
Rwpos63_89 in63 sp89 3183.098862
Rwpos63_90 in63 sp90 11140.846016
Rwpos63_91 in63 sp91 11140.846016
Rwpos63_92 in63 sp92 3183.098862
Rwpos63_93 in63 sp93 3183.098862
Rwpos63_94 in63 sp94 3183.098862
Rwpos63_95 in63 sp95 11140.846016
Rwpos63_96 in63 sp96 11140.846016
Rwpos63_97 in63 sp97 3183.098862
Rwpos63_98 in63 sp98 11140.846016
Rwpos63_99 in63 sp99 3183.098862
Rwpos63_100 in63 sp100 3183.098862
Rwpos64_1 in64 sp1 3183.098862
Rwpos64_2 in64 sp2 3183.098862
Rwpos64_3 in64 sp3 3183.098862
Rwpos64_4 in64 sp4 3183.098862
Rwpos64_5 in64 sp5 11140.846016
Rwpos64_6 in64 sp6 3183.098862
Rwpos64_7 in64 sp7 3183.098862
Rwpos64_8 in64 sp8 3183.098862
Rwpos64_9 in64 sp9 11140.846016
Rwpos64_10 in64 sp10 11140.846016
Rwpos64_11 in64 sp11 3183.098862
Rwpos64_12 in64 sp12 11140.846016
Rwpos64_13 in64 sp13 11140.846016
Rwpos64_14 in64 sp14 3183.098862
Rwpos64_15 in64 sp15 11140.846016
Rwpos64_16 in64 sp16 3183.098862
Rwpos64_17 in64 sp17 3183.098862
Rwpos64_18 in64 sp18 11140.846016
Rwpos64_19 in64 sp19 3183.098862
Rwpos64_20 in64 sp20 3183.098862
Rwpos64_21 in64 sp21 3183.098862
Rwpos64_22 in64 sp22 3183.098862
Rwpos64_23 in64 sp23 3183.098862
Rwpos64_24 in64 sp24 3183.098862
Rwpos64_25 in64 sp25 11140.846016
Rwpos64_26 in64 sp26 11140.846016
Rwpos64_27 in64 sp27 11140.846016
Rwpos64_28 in64 sp28 3183.098862
Rwpos64_29 in64 sp29 3183.098862
Rwpos64_30 in64 sp30 11140.846016
Rwpos64_31 in64 sp31 11140.846016
Rwpos64_32 in64 sp32 11140.846016
Rwpos64_33 in64 sp33 11140.846016
Rwpos64_34 in64 sp34 11140.846016
Rwpos64_35 in64 sp35 11140.846016
Rwpos64_36 in64 sp36 11140.846016
Rwpos64_37 in64 sp37 3183.098862
Rwpos64_38 in64 sp38 3183.098862
Rwpos64_39 in64 sp39 3183.098862
Rwpos64_40 in64 sp40 11140.846016
Rwpos64_41 in64 sp41 11140.846016
Rwpos64_42 in64 sp42 3183.098862
Rwpos64_43 in64 sp43 3183.098862
Rwpos64_44 in64 sp44 11140.846016
Rwpos64_45 in64 sp45 3183.098862
Rwpos64_46 in64 sp46 3183.098862
Rwpos64_47 in64 sp47 3183.098862
Rwpos64_48 in64 sp48 11140.846016
Rwpos64_49 in64 sp49 11140.846016
Rwpos64_50 in64 sp50 3183.098862
Rwpos64_51 in64 sp51 3183.098862
Rwpos64_52 in64 sp52 3183.098862
Rwpos64_53 in64 sp53 3183.098862
Rwpos64_54 in64 sp54 11140.846016
Rwpos64_55 in64 sp55 11140.846016
Rwpos64_56 in64 sp56 11140.846016
Rwpos64_57 in64 sp57 11140.846016
Rwpos64_58 in64 sp58 3183.098862
Rwpos64_59 in64 sp59 11140.846016
Rwpos64_60 in64 sp60 11140.846016
Rwpos64_61 in64 sp61 3183.098862
Rwpos64_62 in64 sp62 11140.846016
Rwpos64_63 in64 sp63 11140.846016
Rwpos64_64 in64 sp64 3183.098862
Rwpos64_65 in64 sp65 3183.098862
Rwpos64_66 in64 sp66 3183.098862
Rwpos64_67 in64 sp67 3183.098862
Rwpos64_68 in64 sp68 3183.098862
Rwpos64_69 in64 sp69 3183.098862
Rwpos64_70 in64 sp70 11140.846016
Rwpos64_71 in64 sp71 3183.098862
Rwpos64_72 in64 sp72 3183.098862
Rwpos64_73 in64 sp73 11140.846016
Rwpos64_74 in64 sp74 3183.098862
Rwpos64_75 in64 sp75 3183.098862
Rwpos64_76 in64 sp76 11140.846016
Rwpos64_77 in64 sp77 11140.846016
Rwpos64_78 in64 sp78 11140.846016
Rwpos64_79 in64 sp79 3183.098862
Rwpos64_80 in64 sp80 11140.846016
Rwpos64_81 in64 sp81 3183.098862
Rwpos64_82 in64 sp82 3183.098862
Rwpos64_83 in64 sp83 3183.098862
Rwpos64_84 in64 sp84 3183.098862
Rwpos64_85 in64 sp85 3183.098862
Rwpos64_86 in64 sp86 11140.846016
Rwpos64_87 in64 sp87 11140.846016
Rwpos64_88 in64 sp88 3183.098862
Rwpos64_89 in64 sp89 3183.098862
Rwpos64_90 in64 sp90 11140.846016
Rwpos64_91 in64 sp91 11140.846016
Rwpos64_92 in64 sp92 11140.846016
Rwpos64_93 in64 sp93 11140.846016
Rwpos64_94 in64 sp94 11140.846016
Rwpos64_95 in64 sp95 3183.098862
Rwpos64_96 in64 sp96 3183.098862
Rwpos64_97 in64 sp97 3183.098862
Rwpos64_98 in64 sp98 3183.098862
Rwpos64_99 in64 sp99 11140.846016
Rwpos64_100 in64 sp100 3183.098862
Rwpos65_1 in65 sp1 3183.098862
Rwpos65_2 in65 sp2 11140.846016
Rwpos65_3 in65 sp3 3183.098862
Rwpos65_4 in65 sp4 3183.098862
Rwpos65_5 in65 sp5 3183.098862
Rwpos65_6 in65 sp6 3183.098862
Rwpos65_7 in65 sp7 11140.846016
Rwpos65_8 in65 sp8 3183.098862
Rwpos65_9 in65 sp9 11140.846016
Rwpos65_10 in65 sp10 11140.846016
Rwpos65_11 in65 sp11 3183.098862
Rwpos65_12 in65 sp12 3183.098862
Rwpos65_13 in65 sp13 3183.098862
Rwpos65_14 in65 sp14 3183.098862
Rwpos65_15 in65 sp15 11140.846016
Rwpos65_16 in65 sp16 3183.098862
Rwpos65_17 in65 sp17 3183.098862
Rwpos65_18 in65 sp18 3183.098862
Rwpos65_19 in65 sp19 3183.098862
Rwpos65_20 in65 sp20 3183.098862
Rwpos65_21 in65 sp21 3183.098862
Rwpos65_22 in65 sp22 11140.846016
Rwpos65_23 in65 sp23 11140.846016
Rwpos65_24 in65 sp24 11140.846016
Rwpos65_25 in65 sp25 11140.846016
Rwpos65_26 in65 sp26 11140.846016
Rwpos65_27 in65 sp27 3183.098862
Rwpos65_28 in65 sp28 3183.098862
Rwpos65_29 in65 sp29 3183.098862
Rwpos65_30 in65 sp30 3183.098862
Rwpos65_31 in65 sp31 3183.098862
Rwpos65_32 in65 sp32 11140.846016
Rwpos65_33 in65 sp33 3183.098862
Rwpos65_34 in65 sp34 3183.098862
Rwpos65_35 in65 sp35 11140.846016
Rwpos65_36 in65 sp36 3183.098862
Rwpos65_37 in65 sp37 3183.098862
Rwpos65_38 in65 sp38 3183.098862
Rwpos65_39 in65 sp39 3183.098862
Rwpos65_40 in65 sp40 3183.098862
Rwpos65_41 in65 sp41 11140.846016
Rwpos65_42 in65 sp42 11140.846016
Rwpos65_43 in65 sp43 3183.098862
Rwpos65_44 in65 sp44 11140.846016
Rwpos65_45 in65 sp45 3183.098862
Rwpos65_46 in65 sp46 3183.098862
Rwpos65_47 in65 sp47 3183.098862
Rwpos65_48 in65 sp48 11140.846016
Rwpos65_49 in65 sp49 3183.098862
Rwpos65_50 in65 sp50 11140.846016
Rwpos65_51 in65 sp51 11140.846016
Rwpos65_52 in65 sp52 3183.098862
Rwpos65_53 in65 sp53 3183.098862
Rwpos65_54 in65 sp54 11140.846016
Rwpos65_55 in65 sp55 3183.098862
Rwpos65_56 in65 sp56 11140.846016
Rwpos65_57 in65 sp57 11140.846016
Rwpos65_58 in65 sp58 11140.846016
Rwpos65_59 in65 sp59 11140.846016
Rwpos65_60 in65 sp60 3183.098862
Rwpos65_61 in65 sp61 11140.846016
Rwpos65_62 in65 sp62 3183.098862
Rwpos65_63 in65 sp63 3183.098862
Rwpos65_64 in65 sp64 11140.846016
Rwpos65_65 in65 sp65 3183.098862
Rwpos65_66 in65 sp66 11140.846016
Rwpos65_67 in65 sp67 3183.098862
Rwpos65_68 in65 sp68 3183.098862
Rwpos65_69 in65 sp69 3183.098862
Rwpos65_70 in65 sp70 11140.846016
Rwpos65_71 in65 sp71 3183.098862
Rwpos65_72 in65 sp72 3183.098862
Rwpos65_73 in65 sp73 3183.098862
Rwpos65_74 in65 sp74 11140.846016
Rwpos65_75 in65 sp75 11140.846016
Rwpos65_76 in65 sp76 3183.098862
Rwpos65_77 in65 sp77 11140.846016
Rwpos65_78 in65 sp78 11140.846016
Rwpos65_79 in65 sp79 3183.098862
Rwpos65_80 in65 sp80 11140.846016
Rwpos65_81 in65 sp81 3183.098862
Rwpos65_82 in65 sp82 11140.846016
Rwpos65_83 in65 sp83 11140.846016
Rwpos65_84 in65 sp84 3183.098862
Rwpos65_85 in65 sp85 3183.098862
Rwpos65_86 in65 sp86 3183.098862
Rwpos65_87 in65 sp87 11140.846016
Rwpos65_88 in65 sp88 3183.098862
Rwpos65_89 in65 sp89 3183.098862
Rwpos65_90 in65 sp90 11140.846016
Rwpos65_91 in65 sp91 11140.846016
Rwpos65_92 in65 sp92 3183.098862
Rwpos65_93 in65 sp93 3183.098862
Rwpos65_94 in65 sp94 11140.846016
Rwpos65_95 in65 sp95 3183.098862
Rwpos65_96 in65 sp96 3183.098862
Rwpos65_97 in65 sp97 3183.098862
Rwpos65_98 in65 sp98 3183.098862
Rwpos65_99 in65 sp99 11140.846016
Rwpos65_100 in65 sp100 3183.098862
Rwpos66_1 in66 sp1 3183.098862
Rwpos66_2 in66 sp2 3183.098862
Rwpos66_3 in66 sp3 11140.846016
Rwpos66_4 in66 sp4 3183.098862
Rwpos66_5 in66 sp5 3183.098862
Rwpos66_6 in66 sp6 3183.098862
Rwpos66_7 in66 sp7 3183.098862
Rwpos66_8 in66 sp8 3183.098862
Rwpos66_9 in66 sp9 3183.098862
Rwpos66_10 in66 sp10 11140.846016
Rwpos66_11 in66 sp11 3183.098862
Rwpos66_12 in66 sp12 3183.098862
Rwpos66_13 in66 sp13 3183.098862
Rwpos66_14 in66 sp14 3183.098862
Rwpos66_15 in66 sp15 11140.846016
Rwpos66_16 in66 sp16 11140.846016
Rwpos66_17 in66 sp17 3183.098862
Rwpos66_18 in66 sp18 11140.846016
Rwpos66_19 in66 sp19 11140.846016
Rwpos66_20 in66 sp20 11140.846016
Rwpos66_21 in66 sp21 3183.098862
Rwpos66_22 in66 sp22 3183.098862
Rwpos66_23 in66 sp23 3183.098862
Rwpos66_24 in66 sp24 3183.098862
Rwpos66_25 in66 sp25 3183.098862
Rwpos66_26 in66 sp26 11140.846016
Rwpos66_27 in66 sp27 3183.098862
Rwpos66_28 in66 sp28 3183.098862
Rwpos66_29 in66 sp29 11140.846016
Rwpos66_30 in66 sp30 11140.846016
Rwpos66_31 in66 sp31 11140.846016
Rwpos66_32 in66 sp32 3183.098862
Rwpos66_33 in66 sp33 3183.098862
Rwpos66_34 in66 sp34 3183.098862
Rwpos66_35 in66 sp35 3183.098862
Rwpos66_36 in66 sp36 11140.846016
Rwpos66_37 in66 sp37 3183.098862
Rwpos66_38 in66 sp38 11140.846016
Rwpos66_39 in66 sp39 3183.098862
Rwpos66_40 in66 sp40 3183.098862
Rwpos66_41 in66 sp41 11140.846016
Rwpos66_42 in66 sp42 3183.098862
Rwpos66_43 in66 sp43 3183.098862
Rwpos66_44 in66 sp44 11140.846016
Rwpos66_45 in66 sp45 11140.846016
Rwpos66_46 in66 sp46 11140.846016
Rwpos66_47 in66 sp47 3183.098862
Rwpos66_48 in66 sp48 3183.098862
Rwpos66_49 in66 sp49 3183.098862
Rwpos66_50 in66 sp50 11140.846016
Rwpos66_51 in66 sp51 3183.098862
Rwpos66_52 in66 sp52 11140.846016
Rwpos66_53 in66 sp53 3183.098862
Rwpos66_54 in66 sp54 3183.098862
Rwpos66_55 in66 sp55 11140.846016
Rwpos66_56 in66 sp56 3183.098862
Rwpos66_57 in66 sp57 3183.098862
Rwpos66_58 in66 sp58 3183.098862
Rwpos66_59 in66 sp59 3183.098862
Rwpos66_60 in66 sp60 3183.098862
Rwpos66_61 in66 sp61 11140.846016
Rwpos66_62 in66 sp62 3183.098862
Rwpos66_63 in66 sp63 11140.846016
Rwpos66_64 in66 sp64 11140.846016
Rwpos66_65 in66 sp65 11140.846016
Rwpos66_66 in66 sp66 11140.846016
Rwpos66_67 in66 sp67 3183.098862
Rwpos66_68 in66 sp68 11140.846016
Rwpos66_69 in66 sp69 3183.098862
Rwpos66_70 in66 sp70 3183.098862
Rwpos66_71 in66 sp71 11140.846016
Rwpos66_72 in66 sp72 3183.098862
Rwpos66_73 in66 sp73 3183.098862
Rwpos66_74 in66 sp74 3183.098862
Rwpos66_75 in66 sp75 3183.098862
Rwpos66_76 in66 sp76 3183.098862
Rwpos66_77 in66 sp77 11140.846016
Rwpos66_78 in66 sp78 11140.846016
Rwpos66_79 in66 sp79 3183.098862
Rwpos66_80 in66 sp80 11140.846016
Rwpos66_81 in66 sp81 3183.098862
Rwpos66_82 in66 sp82 11140.846016
Rwpos66_83 in66 sp83 3183.098862
Rwpos66_84 in66 sp84 11140.846016
Rwpos66_85 in66 sp85 3183.098862
Rwpos66_86 in66 sp86 11140.846016
Rwpos66_87 in66 sp87 11140.846016
Rwpos66_88 in66 sp88 3183.098862
Rwpos66_89 in66 sp89 11140.846016
Rwpos66_90 in66 sp90 3183.098862
Rwpos66_91 in66 sp91 3183.098862
Rwpos66_92 in66 sp92 11140.846016
Rwpos66_93 in66 sp93 11140.846016
Rwpos66_94 in66 sp94 11140.846016
Rwpos66_95 in66 sp95 3183.098862
Rwpos66_96 in66 sp96 11140.846016
Rwpos66_97 in66 sp97 3183.098862
Rwpos66_98 in66 sp98 11140.846016
Rwpos66_99 in66 sp99 3183.098862
Rwpos66_100 in66 sp100 11140.846016
Rwpos67_1 in67 sp1 11140.846016
Rwpos67_2 in67 sp2 11140.846016
Rwpos67_3 in67 sp3 11140.846016
Rwpos67_4 in67 sp4 3183.098862
Rwpos67_5 in67 sp5 3183.098862
Rwpos67_6 in67 sp6 3183.098862
Rwpos67_7 in67 sp7 11140.846016
Rwpos67_8 in67 sp8 3183.098862
Rwpos67_9 in67 sp9 11140.846016
Rwpos67_10 in67 sp10 3183.098862
Rwpos67_11 in67 sp11 11140.846016
Rwpos67_12 in67 sp12 3183.098862
Rwpos67_13 in67 sp13 3183.098862
Rwpos67_14 in67 sp14 11140.846016
Rwpos67_15 in67 sp15 3183.098862
Rwpos67_16 in67 sp16 3183.098862
Rwpos67_17 in67 sp17 3183.098862
Rwpos67_18 in67 sp18 11140.846016
Rwpos67_19 in67 sp19 3183.098862
Rwpos67_20 in67 sp20 11140.846016
Rwpos67_21 in67 sp21 3183.098862
Rwpos67_22 in67 sp22 3183.098862
Rwpos67_23 in67 sp23 11140.846016
Rwpos67_24 in67 sp24 3183.098862
Rwpos67_25 in67 sp25 3183.098862
Rwpos67_26 in67 sp26 3183.098862
Rwpos67_27 in67 sp27 3183.098862
Rwpos67_28 in67 sp28 11140.846016
Rwpos67_29 in67 sp29 3183.098862
Rwpos67_30 in67 sp30 11140.846016
Rwpos67_31 in67 sp31 3183.098862
Rwpos67_32 in67 sp32 3183.098862
Rwpos67_33 in67 sp33 3183.098862
Rwpos67_34 in67 sp34 11140.846016
Rwpos67_35 in67 sp35 3183.098862
Rwpos67_36 in67 sp36 3183.098862
Rwpos67_37 in67 sp37 3183.098862
Rwpos67_38 in67 sp38 3183.098862
Rwpos67_39 in67 sp39 11140.846016
Rwpos67_40 in67 sp40 3183.098862
Rwpos67_41 in67 sp41 3183.098862
Rwpos67_42 in67 sp42 3183.098862
Rwpos67_43 in67 sp43 3183.098862
Rwpos67_44 in67 sp44 3183.098862
Rwpos67_45 in67 sp45 11140.846016
Rwpos67_46 in67 sp46 11140.846016
Rwpos67_47 in67 sp47 11140.846016
Rwpos67_48 in67 sp48 3183.098862
Rwpos67_49 in67 sp49 3183.098862
Rwpos67_50 in67 sp50 11140.846016
Rwpos67_51 in67 sp51 3183.098862
Rwpos67_52 in67 sp52 3183.098862
Rwpos67_53 in67 sp53 3183.098862
Rwpos67_54 in67 sp54 3183.098862
Rwpos67_55 in67 sp55 11140.846016
Rwpos67_56 in67 sp56 11140.846016
Rwpos67_57 in67 sp57 11140.846016
Rwpos67_58 in67 sp58 3183.098862
Rwpos67_59 in67 sp59 11140.846016
Rwpos67_60 in67 sp60 11140.846016
Rwpos67_61 in67 sp61 11140.846016
Rwpos67_62 in67 sp62 11140.846016
Rwpos67_63 in67 sp63 11140.846016
Rwpos67_64 in67 sp64 3183.098862
Rwpos67_65 in67 sp65 11140.846016
Rwpos67_66 in67 sp66 3183.098862
Rwpos67_67 in67 sp67 3183.098862
Rwpos67_68 in67 sp68 3183.098862
Rwpos67_69 in67 sp69 11140.846016
Rwpos67_70 in67 sp70 3183.098862
Rwpos67_71 in67 sp71 11140.846016
Rwpos67_72 in67 sp72 3183.098862
Rwpos67_73 in67 sp73 11140.846016
Rwpos67_74 in67 sp74 3183.098862
Rwpos67_75 in67 sp75 3183.098862
Rwpos67_76 in67 sp76 3183.098862
Rwpos67_77 in67 sp77 11140.846016
Rwpos67_78 in67 sp78 3183.098862
Rwpos67_79 in67 sp79 11140.846016
Rwpos67_80 in67 sp80 3183.098862
Rwpos67_81 in67 sp81 3183.098862
Rwpos67_82 in67 sp82 11140.846016
Rwpos67_83 in67 sp83 11140.846016
Rwpos67_84 in67 sp84 3183.098862
Rwpos67_85 in67 sp85 3183.098862
Rwpos67_86 in67 sp86 11140.846016
Rwpos67_87 in67 sp87 3183.098862
Rwpos67_88 in67 sp88 11140.846016
Rwpos67_89 in67 sp89 11140.846016
Rwpos67_90 in67 sp90 11140.846016
Rwpos67_91 in67 sp91 3183.098862
Rwpos67_92 in67 sp92 3183.098862
Rwpos67_93 in67 sp93 11140.846016
Rwpos67_94 in67 sp94 3183.098862
Rwpos67_95 in67 sp95 11140.846016
Rwpos67_96 in67 sp96 3183.098862
Rwpos67_97 in67 sp97 3183.098862
Rwpos67_98 in67 sp98 11140.846016
Rwpos67_99 in67 sp99 3183.098862
Rwpos67_100 in67 sp100 3183.098862
Rwpos68_1 in68 sp1 11140.846016
Rwpos68_2 in68 sp2 3183.098862
Rwpos68_3 in68 sp3 3183.098862
Rwpos68_4 in68 sp4 3183.098862
Rwpos68_5 in68 sp5 3183.098862
Rwpos68_6 in68 sp6 11140.846016
Rwpos68_7 in68 sp7 11140.846016
Rwpos68_8 in68 sp8 3183.098862
Rwpos68_9 in68 sp9 11140.846016
Rwpos68_10 in68 sp10 3183.098862
Rwpos68_11 in68 sp11 11140.846016
Rwpos68_12 in68 sp12 11140.846016
Rwpos68_13 in68 sp13 3183.098862
Rwpos68_14 in68 sp14 11140.846016
Rwpos68_15 in68 sp15 3183.098862
Rwpos68_16 in68 sp16 3183.098862
Rwpos68_17 in68 sp17 3183.098862
Rwpos68_18 in68 sp18 3183.098862
Rwpos68_19 in68 sp19 11140.846016
Rwpos68_20 in68 sp20 11140.846016
Rwpos68_21 in68 sp21 11140.846016
Rwpos68_22 in68 sp22 3183.098862
Rwpos68_23 in68 sp23 3183.098862
Rwpos68_24 in68 sp24 11140.846016
Rwpos68_25 in68 sp25 3183.098862
Rwpos68_26 in68 sp26 11140.846016
Rwpos68_27 in68 sp27 11140.846016
Rwpos68_28 in68 sp28 11140.846016
Rwpos68_29 in68 sp29 3183.098862
Rwpos68_30 in68 sp30 3183.098862
Rwpos68_31 in68 sp31 11140.846016
Rwpos68_32 in68 sp32 3183.098862
Rwpos68_33 in68 sp33 3183.098862
Rwpos68_34 in68 sp34 11140.846016
Rwpos68_35 in68 sp35 11140.846016
Rwpos68_36 in68 sp36 3183.098862
Rwpos68_37 in68 sp37 3183.098862
Rwpos68_38 in68 sp38 11140.846016
Rwpos68_39 in68 sp39 3183.098862
Rwpos68_40 in68 sp40 3183.098862
Rwpos68_41 in68 sp41 11140.846016
Rwpos68_42 in68 sp42 3183.098862
Rwpos68_43 in68 sp43 11140.846016
Rwpos68_44 in68 sp44 3183.098862
Rwpos68_45 in68 sp45 3183.098862
Rwpos68_46 in68 sp46 3183.098862
Rwpos68_47 in68 sp47 11140.846016
Rwpos68_48 in68 sp48 3183.098862
Rwpos68_49 in68 sp49 3183.098862
Rwpos68_50 in68 sp50 3183.098862
Rwpos68_51 in68 sp51 11140.846016
Rwpos68_52 in68 sp52 11140.846016
Rwpos68_53 in68 sp53 3183.098862
Rwpos68_54 in68 sp54 3183.098862
Rwpos68_55 in68 sp55 11140.846016
Rwpos68_56 in68 sp56 3183.098862
Rwpos68_57 in68 sp57 3183.098862
Rwpos68_58 in68 sp58 3183.098862
Rwpos68_59 in68 sp59 3183.098862
Rwpos68_60 in68 sp60 11140.846016
Rwpos68_61 in68 sp61 3183.098862
Rwpos68_62 in68 sp62 11140.846016
Rwpos68_63 in68 sp63 11140.846016
Rwpos68_64 in68 sp64 11140.846016
Rwpos68_65 in68 sp65 3183.098862
Rwpos68_66 in68 sp66 11140.846016
Rwpos68_67 in68 sp67 3183.098862
Rwpos68_68 in68 sp68 11140.846016
Rwpos68_69 in68 sp69 11140.846016
Rwpos68_70 in68 sp70 3183.098862
Rwpos68_71 in68 sp71 11140.846016
Rwpos68_72 in68 sp72 3183.098862
Rwpos68_73 in68 sp73 3183.098862
Rwpos68_74 in68 sp74 11140.846016
Rwpos68_75 in68 sp75 11140.846016
Rwpos68_76 in68 sp76 3183.098862
Rwpos68_77 in68 sp77 11140.846016
Rwpos68_78 in68 sp78 11140.846016
Rwpos68_79 in68 sp79 11140.846016
Rwpos68_80 in68 sp80 3183.098862
Rwpos68_81 in68 sp81 3183.098862
Rwpos68_82 in68 sp82 3183.098862
Rwpos68_83 in68 sp83 11140.846016
Rwpos68_84 in68 sp84 3183.098862
Rwpos68_85 in68 sp85 3183.098862
Rwpos68_86 in68 sp86 3183.098862
Rwpos68_87 in68 sp87 3183.098862
Rwpos68_88 in68 sp88 3183.098862
Rwpos68_89 in68 sp89 3183.098862
Rwpos68_90 in68 sp90 11140.846016
Rwpos68_91 in68 sp91 11140.846016
Rwpos68_92 in68 sp92 11140.846016
Rwpos68_93 in68 sp93 11140.846016
Rwpos68_94 in68 sp94 3183.098862
Rwpos68_95 in68 sp95 11140.846016
Rwpos68_96 in68 sp96 3183.098862
Rwpos68_97 in68 sp97 3183.098862
Rwpos68_98 in68 sp98 11140.846016
Rwpos68_99 in68 sp99 11140.846016
Rwpos68_100 in68 sp100 11140.846016
Rwpos69_1 in69 sp1 3183.098862
Rwpos69_2 in69 sp2 3183.098862
Rwpos69_3 in69 sp3 11140.846016
Rwpos69_4 in69 sp4 3183.098862
Rwpos69_5 in69 sp5 3183.098862
Rwpos69_6 in69 sp6 3183.098862
Rwpos69_7 in69 sp7 3183.098862
Rwpos69_8 in69 sp8 3183.098862
Rwpos69_9 in69 sp9 11140.846016
Rwpos69_10 in69 sp10 11140.846016
Rwpos69_11 in69 sp11 3183.098862
Rwpos69_12 in69 sp12 11140.846016
Rwpos69_13 in69 sp13 3183.098862
Rwpos69_14 in69 sp14 3183.098862
Rwpos69_15 in69 sp15 3183.098862
Rwpos69_16 in69 sp16 3183.098862
Rwpos69_17 in69 sp17 3183.098862
Rwpos69_18 in69 sp18 11140.846016
Rwpos69_19 in69 sp19 3183.098862
Rwpos69_20 in69 sp20 3183.098862
Rwpos69_21 in69 sp21 11140.846016
Rwpos69_22 in69 sp22 3183.098862
Rwpos69_23 in69 sp23 3183.098862
Rwpos69_24 in69 sp24 11140.846016
Rwpos69_25 in69 sp25 11140.846016
Rwpos69_26 in69 sp26 11140.846016
Rwpos69_27 in69 sp27 3183.098862
Rwpos69_28 in69 sp28 11140.846016
Rwpos69_29 in69 sp29 3183.098862
Rwpos69_30 in69 sp30 3183.098862
Rwpos69_31 in69 sp31 3183.098862
Rwpos69_32 in69 sp32 3183.098862
Rwpos69_33 in69 sp33 3183.098862
Rwpos69_34 in69 sp34 11140.846016
Rwpos69_35 in69 sp35 11140.846016
Rwpos69_36 in69 sp36 3183.098862
Rwpos69_37 in69 sp37 3183.098862
Rwpos69_38 in69 sp38 3183.098862
Rwpos69_39 in69 sp39 3183.098862
Rwpos69_40 in69 sp40 11140.846016
Rwpos69_41 in69 sp41 11140.846016
Rwpos69_42 in69 sp42 11140.846016
Rwpos69_43 in69 sp43 3183.098862
Rwpos69_44 in69 sp44 11140.846016
Rwpos69_45 in69 sp45 3183.098862
Rwpos69_46 in69 sp46 3183.098862
Rwpos69_47 in69 sp47 3183.098862
Rwpos69_48 in69 sp48 3183.098862
Rwpos69_49 in69 sp49 3183.098862
Rwpos69_50 in69 sp50 11140.846016
Rwpos69_51 in69 sp51 3183.098862
Rwpos69_52 in69 sp52 3183.098862
Rwpos69_53 in69 sp53 3183.098862
Rwpos69_54 in69 sp54 11140.846016
Rwpos69_55 in69 sp55 11140.846016
Rwpos69_56 in69 sp56 11140.846016
Rwpos69_57 in69 sp57 3183.098862
Rwpos69_58 in69 sp58 11140.846016
Rwpos69_59 in69 sp59 11140.846016
Rwpos69_60 in69 sp60 11140.846016
Rwpos69_61 in69 sp61 3183.098862
Rwpos69_62 in69 sp62 3183.098862
Rwpos69_63 in69 sp63 3183.098862
Rwpos69_64 in69 sp64 3183.098862
Rwpos69_65 in69 sp65 3183.098862
Rwpos69_66 in69 sp66 3183.098862
Rwpos69_67 in69 sp67 11140.846016
Rwpos69_68 in69 sp68 3183.098862
Rwpos69_69 in69 sp69 3183.098862
Rwpos69_70 in69 sp70 3183.098862
Rwpos69_71 in69 sp71 3183.098862
Rwpos69_72 in69 sp72 11140.846016
Rwpos69_73 in69 sp73 11140.846016
Rwpos69_74 in69 sp74 11140.846016
Rwpos69_75 in69 sp75 11140.846016
Rwpos69_76 in69 sp76 11140.846016
Rwpos69_77 in69 sp77 11140.846016
Rwpos69_78 in69 sp78 3183.098862
Rwpos69_79 in69 sp79 11140.846016
Rwpos69_80 in69 sp80 11140.846016
Rwpos69_81 in69 sp81 3183.098862
Rwpos69_82 in69 sp82 11140.846016
Rwpos69_83 in69 sp83 11140.846016
Rwpos69_84 in69 sp84 3183.098862
Rwpos69_85 in69 sp85 3183.098862
Rwpos69_86 in69 sp86 11140.846016
Rwpos69_87 in69 sp87 11140.846016
Rwpos69_88 in69 sp88 3183.098862
Rwpos69_89 in69 sp89 11140.846016
Rwpos69_90 in69 sp90 11140.846016
Rwpos69_91 in69 sp91 3183.098862
Rwpos69_92 in69 sp92 11140.846016
Rwpos69_93 in69 sp93 3183.098862
Rwpos69_94 in69 sp94 3183.098862
Rwpos69_95 in69 sp95 3183.098862
Rwpos69_96 in69 sp96 11140.846016
Rwpos69_97 in69 sp97 11140.846016
Rwpos69_98 in69 sp98 11140.846016
Rwpos69_99 in69 sp99 11140.846016
Rwpos69_100 in69 sp100 3183.098862
Rwpos70_1 in70 sp1 3183.098862
Rwpos70_2 in70 sp2 3183.098862
Rwpos70_3 in70 sp3 3183.098862
Rwpos70_4 in70 sp4 11140.846016
Rwpos70_5 in70 sp5 11140.846016
Rwpos70_6 in70 sp6 11140.846016
Rwpos70_7 in70 sp7 11140.846016
Rwpos70_8 in70 sp8 11140.846016
Rwpos70_9 in70 sp9 11140.846016
Rwpos70_10 in70 sp10 3183.098862
Rwpos70_11 in70 sp11 3183.098862
Rwpos70_12 in70 sp12 11140.846016
Rwpos70_13 in70 sp13 3183.098862
Rwpos70_14 in70 sp14 11140.846016
Rwpos70_15 in70 sp15 11140.846016
Rwpos70_16 in70 sp16 3183.098862
Rwpos70_17 in70 sp17 3183.098862
Rwpos70_18 in70 sp18 11140.846016
Rwpos70_19 in70 sp19 11140.846016
Rwpos70_20 in70 sp20 3183.098862
Rwpos70_21 in70 sp21 3183.098862
Rwpos70_22 in70 sp22 11140.846016
Rwpos70_23 in70 sp23 3183.098862
Rwpos70_24 in70 sp24 3183.098862
Rwpos70_25 in70 sp25 11140.846016
Rwpos70_26 in70 sp26 11140.846016
Rwpos70_27 in70 sp27 3183.098862
Rwpos70_28 in70 sp28 11140.846016
Rwpos70_29 in70 sp29 3183.098862
Rwpos70_30 in70 sp30 11140.846016
Rwpos70_31 in70 sp31 11140.846016
Rwpos70_32 in70 sp32 11140.846016
Rwpos70_33 in70 sp33 3183.098862
Rwpos70_34 in70 sp34 3183.098862
Rwpos70_35 in70 sp35 11140.846016
Rwpos70_36 in70 sp36 11140.846016
Rwpos70_37 in70 sp37 3183.098862
Rwpos70_38 in70 sp38 3183.098862
Rwpos70_39 in70 sp39 11140.846016
Rwpos70_40 in70 sp40 3183.098862
Rwpos70_41 in70 sp41 11140.846016
Rwpos70_42 in70 sp42 11140.846016
Rwpos70_43 in70 sp43 3183.098862
Rwpos70_44 in70 sp44 11140.846016
Rwpos70_45 in70 sp45 3183.098862
Rwpos70_46 in70 sp46 11140.846016
Rwpos70_47 in70 sp47 3183.098862
Rwpos70_48 in70 sp48 11140.846016
Rwpos70_49 in70 sp49 3183.098862
Rwpos70_50 in70 sp50 11140.846016
Rwpos70_51 in70 sp51 3183.098862
Rwpos70_52 in70 sp52 3183.098862
Rwpos70_53 in70 sp53 3183.098862
Rwpos70_54 in70 sp54 11140.846016
Rwpos70_55 in70 sp55 11140.846016
Rwpos70_56 in70 sp56 3183.098862
Rwpos70_57 in70 sp57 3183.098862
Rwpos70_58 in70 sp58 11140.846016
Rwpos70_59 in70 sp59 3183.098862
Rwpos70_60 in70 sp60 11140.846016
Rwpos70_61 in70 sp61 11140.846016
Rwpos70_62 in70 sp62 11140.846016
Rwpos70_63 in70 sp63 11140.846016
Rwpos70_64 in70 sp64 3183.098862
Rwpos70_65 in70 sp65 3183.098862
Rwpos70_66 in70 sp66 11140.846016
Rwpos70_67 in70 sp67 11140.846016
Rwpos70_68 in70 sp68 11140.846016
Rwpos70_69 in70 sp69 3183.098862
Rwpos70_70 in70 sp70 11140.846016
Rwpos70_71 in70 sp71 3183.098862
Rwpos70_72 in70 sp72 3183.098862
Rwpos70_73 in70 sp73 3183.098862
Rwpos70_74 in70 sp74 11140.846016
Rwpos70_75 in70 sp75 3183.098862
Rwpos70_76 in70 sp76 3183.098862
Rwpos70_77 in70 sp77 11140.846016
Rwpos70_78 in70 sp78 11140.846016
Rwpos70_79 in70 sp79 11140.846016
Rwpos70_80 in70 sp80 3183.098862
Rwpos70_81 in70 sp81 11140.846016
Rwpos70_82 in70 sp82 11140.846016
Rwpos70_83 in70 sp83 3183.098862
Rwpos70_84 in70 sp84 11140.846016
Rwpos70_85 in70 sp85 3183.098862
Rwpos70_86 in70 sp86 11140.846016
Rwpos70_87 in70 sp87 11140.846016
Rwpos70_88 in70 sp88 3183.098862
Rwpos70_89 in70 sp89 3183.098862
Rwpos70_90 in70 sp90 11140.846016
Rwpos70_91 in70 sp91 3183.098862
Rwpos70_92 in70 sp92 11140.846016
Rwpos70_93 in70 sp93 11140.846016
Rwpos70_94 in70 sp94 3183.098862
Rwpos70_95 in70 sp95 11140.846016
Rwpos70_96 in70 sp96 3183.098862
Rwpos70_97 in70 sp97 3183.098862
Rwpos70_98 in70 sp98 11140.846016
Rwpos70_99 in70 sp99 3183.098862
Rwpos70_100 in70 sp100 11140.846016
Rwpos71_1 in71 sp1 3183.098862
Rwpos71_2 in71 sp2 11140.846016
Rwpos71_3 in71 sp3 3183.098862
Rwpos71_4 in71 sp4 3183.098862
Rwpos71_5 in71 sp5 3183.098862
Rwpos71_6 in71 sp6 3183.098862
Rwpos71_7 in71 sp7 11140.846016
Rwpos71_8 in71 sp8 3183.098862
Rwpos71_9 in71 sp9 11140.846016
Rwpos71_10 in71 sp10 11140.846016
Rwpos71_11 in71 sp11 3183.098862
Rwpos71_12 in71 sp12 11140.846016
Rwpos71_13 in71 sp13 3183.098862
Rwpos71_14 in71 sp14 11140.846016
Rwpos71_15 in71 sp15 11140.846016
Rwpos71_16 in71 sp16 11140.846016
Rwpos71_17 in71 sp17 3183.098862
Rwpos71_18 in71 sp18 3183.098862
Rwpos71_19 in71 sp19 3183.098862
Rwpos71_20 in71 sp20 11140.846016
Rwpos71_21 in71 sp21 3183.098862
Rwpos71_22 in71 sp22 3183.098862
Rwpos71_23 in71 sp23 3183.098862
Rwpos71_24 in71 sp24 3183.098862
Rwpos71_25 in71 sp25 11140.846016
Rwpos71_26 in71 sp26 3183.098862
Rwpos71_27 in71 sp27 11140.846016
Rwpos71_28 in71 sp28 11140.846016
Rwpos71_29 in71 sp29 3183.098862
Rwpos71_30 in71 sp30 11140.846016
Rwpos71_31 in71 sp31 3183.098862
Rwpos71_32 in71 sp32 11140.846016
Rwpos71_33 in71 sp33 3183.098862
Rwpos71_34 in71 sp34 11140.846016
Rwpos71_35 in71 sp35 3183.098862
Rwpos71_36 in71 sp36 11140.846016
Rwpos71_37 in71 sp37 3183.098862
Rwpos71_38 in71 sp38 3183.098862
Rwpos71_39 in71 sp39 11140.846016
Rwpos71_40 in71 sp40 11140.846016
Rwpos71_41 in71 sp41 11140.846016
Rwpos71_42 in71 sp42 11140.846016
Rwpos71_43 in71 sp43 3183.098862
Rwpos71_44 in71 sp44 11140.846016
Rwpos71_45 in71 sp45 3183.098862
Rwpos71_46 in71 sp46 11140.846016
Rwpos71_47 in71 sp47 3183.098862
Rwpos71_48 in71 sp48 11140.846016
Rwpos71_49 in71 sp49 3183.098862
Rwpos71_50 in71 sp50 11140.846016
Rwpos71_51 in71 sp51 3183.098862
Rwpos71_52 in71 sp52 3183.098862
Rwpos71_53 in71 sp53 3183.098862
Rwpos71_54 in71 sp54 3183.098862
Rwpos71_55 in71 sp55 3183.098862
Rwpos71_56 in71 sp56 3183.098862
Rwpos71_57 in71 sp57 11140.846016
Rwpos71_58 in71 sp58 3183.098862
Rwpos71_59 in71 sp59 3183.098862
Rwpos71_60 in71 sp60 3183.098862
Rwpos71_61 in71 sp61 11140.846016
Rwpos71_62 in71 sp62 11140.846016
Rwpos71_63 in71 sp63 11140.846016
Rwpos71_64 in71 sp64 3183.098862
Rwpos71_65 in71 sp65 11140.846016
Rwpos71_66 in71 sp66 11140.846016
Rwpos71_67 in71 sp67 3183.098862
Rwpos71_68 in71 sp68 3183.098862
Rwpos71_69 in71 sp69 3183.098862
Rwpos71_70 in71 sp70 3183.098862
Rwpos71_71 in71 sp71 11140.846016
Rwpos71_72 in71 sp72 11140.846016
Rwpos71_73 in71 sp73 11140.846016
Rwpos71_74 in71 sp74 11140.846016
Rwpos71_75 in71 sp75 3183.098862
Rwpos71_76 in71 sp76 11140.846016
Rwpos71_77 in71 sp77 11140.846016
Rwpos71_78 in71 sp78 11140.846016
Rwpos71_79 in71 sp79 3183.098862
Rwpos71_80 in71 sp80 3183.098862
Rwpos71_81 in71 sp81 11140.846016
Rwpos71_82 in71 sp82 11140.846016
Rwpos71_83 in71 sp83 3183.098862
Rwpos71_84 in71 sp84 11140.846016
Rwpos71_85 in71 sp85 3183.098862
Rwpos71_86 in71 sp86 3183.098862
Rwpos71_87 in71 sp87 11140.846016
Rwpos71_88 in71 sp88 3183.098862
Rwpos71_89 in71 sp89 3183.098862
Rwpos71_90 in71 sp90 11140.846016
Rwpos71_91 in71 sp91 3183.098862
Rwpos71_92 in71 sp92 11140.846016
Rwpos71_93 in71 sp93 11140.846016
Rwpos71_94 in71 sp94 11140.846016
Rwpos71_95 in71 sp95 3183.098862
Rwpos71_96 in71 sp96 3183.098862
Rwpos71_97 in71 sp97 11140.846016
Rwpos71_98 in71 sp98 11140.846016
Rwpos71_99 in71 sp99 3183.098862
Rwpos71_100 in71 sp100 11140.846016
Rwpos72_1 in72 sp1 3183.098862
Rwpos72_2 in72 sp2 3183.098862
Rwpos72_3 in72 sp3 11140.846016
Rwpos72_4 in72 sp4 11140.846016
Rwpos72_5 in72 sp5 3183.098862
Rwpos72_6 in72 sp6 3183.098862
Rwpos72_7 in72 sp7 3183.098862
Rwpos72_8 in72 sp8 3183.098862
Rwpos72_9 in72 sp9 3183.098862
Rwpos72_10 in72 sp10 11140.846016
Rwpos72_11 in72 sp11 11140.846016
Rwpos72_12 in72 sp12 11140.846016
Rwpos72_13 in72 sp13 3183.098862
Rwpos72_14 in72 sp14 11140.846016
Rwpos72_15 in72 sp15 3183.098862
Rwpos72_16 in72 sp16 3183.098862
Rwpos72_17 in72 sp17 3183.098862
Rwpos72_18 in72 sp18 3183.098862
Rwpos72_19 in72 sp19 11140.846016
Rwpos72_20 in72 sp20 11140.846016
Rwpos72_21 in72 sp21 3183.098862
Rwpos72_22 in72 sp22 3183.098862
Rwpos72_23 in72 sp23 3183.098862
Rwpos72_24 in72 sp24 3183.098862
Rwpos72_25 in72 sp25 3183.098862
Rwpos72_26 in72 sp26 11140.846016
Rwpos72_27 in72 sp27 11140.846016
Rwpos72_28 in72 sp28 3183.098862
Rwpos72_29 in72 sp29 11140.846016
Rwpos72_30 in72 sp30 11140.846016
Rwpos72_31 in72 sp31 3183.098862
Rwpos72_32 in72 sp32 11140.846016
Rwpos72_33 in72 sp33 11140.846016
Rwpos72_34 in72 sp34 3183.098862
Rwpos72_35 in72 sp35 3183.098862
Rwpos72_36 in72 sp36 11140.846016
Rwpos72_37 in72 sp37 11140.846016
Rwpos72_38 in72 sp38 11140.846016
Rwpos72_39 in72 sp39 3183.098862
Rwpos72_40 in72 sp40 11140.846016
Rwpos72_41 in72 sp41 11140.846016
Rwpos72_42 in72 sp42 3183.098862
Rwpos72_43 in72 sp43 3183.098862
Rwpos72_44 in72 sp44 3183.098862
Rwpos72_45 in72 sp45 3183.098862
Rwpos72_46 in72 sp46 11140.846016
Rwpos72_47 in72 sp47 11140.846016
Rwpos72_48 in72 sp48 11140.846016
Rwpos72_49 in72 sp49 3183.098862
Rwpos72_50 in72 sp50 3183.098862
Rwpos72_51 in72 sp51 11140.846016
Rwpos72_52 in72 sp52 3183.098862
Rwpos72_53 in72 sp53 11140.846016
Rwpos72_54 in72 sp54 11140.846016
Rwpos72_55 in72 sp55 3183.098862
Rwpos72_56 in72 sp56 3183.098862
Rwpos72_57 in72 sp57 11140.846016
Rwpos72_58 in72 sp58 3183.098862
Rwpos72_59 in72 sp59 3183.098862
Rwpos72_60 in72 sp60 3183.098862
Rwpos72_61 in72 sp61 11140.846016
Rwpos72_62 in72 sp62 11140.846016
Rwpos72_63 in72 sp63 3183.098862
Rwpos72_64 in72 sp64 3183.098862
Rwpos72_65 in72 sp65 11140.846016
Rwpos72_66 in72 sp66 3183.098862
Rwpos72_67 in72 sp67 3183.098862
Rwpos72_68 in72 sp68 3183.098862
Rwpos72_69 in72 sp69 11140.846016
Rwpos72_70 in72 sp70 11140.846016
Rwpos72_71 in72 sp71 11140.846016
Rwpos72_72 in72 sp72 11140.846016
Rwpos72_73 in72 sp73 3183.098862
Rwpos72_74 in72 sp74 11140.846016
Rwpos72_75 in72 sp75 3183.098862
Rwpos72_76 in72 sp76 3183.098862
Rwpos72_77 in72 sp77 11140.846016
Rwpos72_78 in72 sp78 3183.098862
Rwpos72_79 in72 sp79 11140.846016
Rwpos72_80 in72 sp80 11140.846016
Rwpos72_81 in72 sp81 11140.846016
Rwpos72_82 in72 sp82 11140.846016
Rwpos72_83 in72 sp83 11140.846016
Rwpos72_84 in72 sp84 11140.846016
Rwpos72_85 in72 sp85 3183.098862
Rwpos72_86 in72 sp86 11140.846016
Rwpos72_87 in72 sp87 3183.098862
Rwpos72_88 in72 sp88 3183.098862
Rwpos72_89 in72 sp89 3183.098862
Rwpos72_90 in72 sp90 11140.846016
Rwpos72_91 in72 sp91 11140.846016
Rwpos72_92 in72 sp92 11140.846016
Rwpos72_93 in72 sp93 11140.846016
Rwpos72_94 in72 sp94 11140.846016
Rwpos72_95 in72 sp95 3183.098862
Rwpos72_96 in72 sp96 11140.846016
Rwpos72_97 in72 sp97 11140.846016
Rwpos72_98 in72 sp98 3183.098862
Rwpos72_99 in72 sp99 3183.098862
Rwpos72_100 in72 sp100 11140.846016
Rwpos73_1 in73 sp1 11140.846016
Rwpos73_2 in73 sp2 3183.098862
Rwpos73_3 in73 sp3 3183.098862
Rwpos73_4 in73 sp4 11140.846016
Rwpos73_5 in73 sp5 3183.098862
Rwpos73_6 in73 sp6 11140.846016
Rwpos73_7 in73 sp7 11140.846016
Rwpos73_8 in73 sp8 3183.098862
Rwpos73_9 in73 sp9 3183.098862
Rwpos73_10 in73 sp10 3183.098862
Rwpos73_11 in73 sp11 3183.098862
Rwpos73_12 in73 sp12 3183.098862
Rwpos73_13 in73 sp13 3183.098862
Rwpos73_14 in73 sp14 3183.098862
Rwpos73_15 in73 sp15 3183.098862
Rwpos73_16 in73 sp16 3183.098862
Rwpos73_17 in73 sp17 11140.846016
Rwpos73_18 in73 sp18 11140.846016
Rwpos73_19 in73 sp19 3183.098862
Rwpos73_20 in73 sp20 11140.846016
Rwpos73_21 in73 sp21 11140.846016
Rwpos73_22 in73 sp22 3183.098862
Rwpos73_23 in73 sp23 3183.098862
Rwpos73_24 in73 sp24 11140.846016
Rwpos73_25 in73 sp25 11140.846016
Rwpos73_26 in73 sp26 11140.846016
Rwpos73_27 in73 sp27 3183.098862
Rwpos73_28 in73 sp28 3183.098862
Rwpos73_29 in73 sp29 11140.846016
Rwpos73_30 in73 sp30 11140.846016
Rwpos73_31 in73 sp31 3183.098862
Rwpos73_32 in73 sp32 3183.098862
Rwpos73_33 in73 sp33 11140.846016
Rwpos73_34 in73 sp34 11140.846016
Rwpos73_35 in73 sp35 3183.098862
Rwpos73_36 in73 sp36 11140.846016
Rwpos73_37 in73 sp37 3183.098862
Rwpos73_38 in73 sp38 3183.098862
Rwpos73_39 in73 sp39 11140.846016
Rwpos73_40 in73 sp40 11140.846016
Rwpos73_41 in73 sp41 11140.846016
Rwpos73_42 in73 sp42 11140.846016
Rwpos73_43 in73 sp43 11140.846016
Rwpos73_44 in73 sp44 3183.098862
Rwpos73_45 in73 sp45 3183.098862
Rwpos73_46 in73 sp46 11140.846016
Rwpos73_47 in73 sp47 11140.846016
Rwpos73_48 in73 sp48 3183.098862
Rwpos73_49 in73 sp49 11140.846016
Rwpos73_50 in73 sp50 11140.846016
Rwpos73_51 in73 sp51 11140.846016
Rwpos73_52 in73 sp52 3183.098862
Rwpos73_53 in73 sp53 3183.098862
Rwpos73_54 in73 sp54 3183.098862
Rwpos73_55 in73 sp55 3183.098862
Rwpos73_56 in73 sp56 3183.098862
Rwpos73_57 in73 sp57 3183.098862
Rwpos73_58 in73 sp58 3183.098862
Rwpos73_59 in73 sp59 3183.098862
Rwpos73_60 in73 sp60 11140.846016
Rwpos73_61 in73 sp61 3183.098862
Rwpos73_62 in73 sp62 3183.098862
Rwpos73_63 in73 sp63 3183.098862
Rwpos73_64 in73 sp64 3183.098862
Rwpos73_65 in73 sp65 3183.098862
Rwpos73_66 in73 sp66 11140.846016
Rwpos73_67 in73 sp67 3183.098862
Rwpos73_68 in73 sp68 3183.098862
Rwpos73_69 in73 sp69 3183.098862
Rwpos73_70 in73 sp70 3183.098862
Rwpos73_71 in73 sp71 11140.846016
Rwpos73_72 in73 sp72 11140.846016
Rwpos73_73 in73 sp73 3183.098862
Rwpos73_74 in73 sp74 11140.846016
Rwpos73_75 in73 sp75 11140.846016
Rwpos73_76 in73 sp76 11140.846016
Rwpos73_77 in73 sp77 3183.098862
Rwpos73_78 in73 sp78 3183.098862
Rwpos73_79 in73 sp79 11140.846016
Rwpos73_80 in73 sp80 11140.846016
Rwpos73_81 in73 sp81 3183.098862
Rwpos73_82 in73 sp82 3183.098862
Rwpos73_83 in73 sp83 3183.098862
Rwpos73_84 in73 sp84 3183.098862
Rwpos73_85 in73 sp85 11140.846016
Rwpos73_86 in73 sp86 3183.098862
Rwpos73_87 in73 sp87 3183.098862
Rwpos73_88 in73 sp88 3183.098862
Rwpos73_89 in73 sp89 11140.846016
Rwpos73_90 in73 sp90 3183.098862
Rwpos73_91 in73 sp91 3183.098862
Rwpos73_92 in73 sp92 11140.846016
Rwpos73_93 in73 sp93 3183.098862
Rwpos73_94 in73 sp94 3183.098862
Rwpos73_95 in73 sp95 11140.846016
Rwpos73_96 in73 sp96 11140.846016
Rwpos73_97 in73 sp97 3183.098862
Rwpos73_98 in73 sp98 11140.846016
Rwpos73_99 in73 sp99 3183.098862
Rwpos73_100 in73 sp100 3183.098862
Rwpos74_1 in74 sp1 3183.098862
Rwpos74_2 in74 sp2 3183.098862
Rwpos74_3 in74 sp3 3183.098862
Rwpos74_4 in74 sp4 11140.846016
Rwpos74_5 in74 sp5 3183.098862
Rwpos74_6 in74 sp6 11140.846016
Rwpos74_7 in74 sp7 3183.098862
Rwpos74_8 in74 sp8 11140.846016
Rwpos74_9 in74 sp9 3183.098862
Rwpos74_10 in74 sp10 3183.098862
Rwpos74_11 in74 sp11 3183.098862
Rwpos74_12 in74 sp12 11140.846016
Rwpos74_13 in74 sp13 3183.098862
Rwpos74_14 in74 sp14 11140.846016
Rwpos74_15 in74 sp15 11140.846016
Rwpos74_16 in74 sp16 3183.098862
Rwpos74_17 in74 sp17 3183.098862
Rwpos74_18 in74 sp18 11140.846016
Rwpos74_19 in74 sp19 3183.098862
Rwpos74_20 in74 sp20 3183.098862
Rwpos74_21 in74 sp21 11140.846016
Rwpos74_22 in74 sp22 3183.098862
Rwpos74_23 in74 sp23 3183.098862
Rwpos74_24 in74 sp24 11140.846016
Rwpos74_25 in74 sp25 3183.098862
Rwpos74_26 in74 sp26 3183.098862
Rwpos74_27 in74 sp27 11140.846016
Rwpos74_28 in74 sp28 11140.846016
Rwpos74_29 in74 sp29 3183.098862
Rwpos74_30 in74 sp30 11140.846016
Rwpos74_31 in74 sp31 11140.846016
Rwpos74_32 in74 sp32 3183.098862
Rwpos74_33 in74 sp33 3183.098862
Rwpos74_34 in74 sp34 3183.098862
Rwpos74_35 in74 sp35 3183.098862
Rwpos74_36 in74 sp36 11140.846016
Rwpos74_37 in74 sp37 3183.098862
Rwpos74_38 in74 sp38 3183.098862
Rwpos74_39 in74 sp39 3183.098862
Rwpos74_40 in74 sp40 11140.846016
Rwpos74_41 in74 sp41 3183.098862
Rwpos74_42 in74 sp42 3183.098862
Rwpos74_43 in74 sp43 3183.098862
Rwpos74_44 in74 sp44 11140.846016
Rwpos74_45 in74 sp45 3183.098862
Rwpos74_46 in74 sp46 11140.846016
Rwpos74_47 in74 sp47 11140.846016
Rwpos74_48 in74 sp48 3183.098862
Rwpos74_49 in74 sp49 3183.098862
Rwpos74_50 in74 sp50 11140.846016
Rwpos74_51 in74 sp51 11140.846016
Rwpos74_52 in74 sp52 11140.846016
Rwpos74_53 in74 sp53 3183.098862
Rwpos74_54 in74 sp54 3183.098862
Rwpos74_55 in74 sp55 3183.098862
Rwpos74_56 in74 sp56 3183.098862
Rwpos74_57 in74 sp57 11140.846016
Rwpos74_58 in74 sp58 11140.846016
Rwpos74_59 in74 sp59 3183.098862
Rwpos74_60 in74 sp60 11140.846016
Rwpos74_61 in74 sp61 3183.098862
Rwpos74_62 in74 sp62 11140.846016
Rwpos74_63 in74 sp63 11140.846016
Rwpos74_64 in74 sp64 11140.846016
Rwpos74_65 in74 sp65 3183.098862
Rwpos74_66 in74 sp66 3183.098862
Rwpos74_67 in74 sp67 3183.098862
Rwpos74_68 in74 sp68 3183.098862
Rwpos74_69 in74 sp69 3183.098862
Rwpos74_70 in74 sp70 11140.846016
Rwpos74_71 in74 sp71 11140.846016
Rwpos74_72 in74 sp72 3183.098862
Rwpos74_73 in74 sp73 3183.098862
Rwpos74_74 in74 sp74 11140.846016
Rwpos74_75 in74 sp75 3183.098862
Rwpos74_76 in74 sp76 11140.846016
Rwpos74_77 in74 sp77 3183.098862
Rwpos74_78 in74 sp78 11140.846016
Rwpos74_79 in74 sp79 3183.098862
Rwpos74_80 in74 sp80 11140.846016
Rwpos74_81 in74 sp81 3183.098862
Rwpos74_82 in74 sp82 3183.098862
Rwpos74_83 in74 sp83 11140.846016
Rwpos74_84 in74 sp84 3183.098862
Rwpos74_85 in74 sp85 3183.098862
Rwpos74_86 in74 sp86 3183.098862
Rwpos74_87 in74 sp87 3183.098862
Rwpos74_88 in74 sp88 3183.098862
Rwpos74_89 in74 sp89 3183.098862
Rwpos74_90 in74 sp90 11140.846016
Rwpos74_91 in74 sp91 3183.098862
Rwpos74_92 in74 sp92 3183.098862
Rwpos74_93 in74 sp93 3183.098862
Rwpos74_94 in74 sp94 11140.846016
Rwpos74_95 in74 sp95 3183.098862
Rwpos74_96 in74 sp96 11140.846016
Rwpos74_97 in74 sp97 11140.846016
Rwpos74_98 in74 sp98 3183.098862
Rwpos74_99 in74 sp99 11140.846016
Rwpos74_100 in74 sp100 11140.846016
Rwpos75_1 in75 sp1 3183.098862
Rwpos75_2 in75 sp2 11140.846016
Rwpos75_3 in75 sp3 3183.098862
Rwpos75_4 in75 sp4 3183.098862
Rwpos75_5 in75 sp5 3183.098862
Rwpos75_6 in75 sp6 11140.846016
Rwpos75_7 in75 sp7 3183.098862
Rwpos75_8 in75 sp8 11140.846016
Rwpos75_9 in75 sp9 11140.846016
Rwpos75_10 in75 sp10 11140.846016
Rwpos75_11 in75 sp11 3183.098862
Rwpos75_12 in75 sp12 3183.098862
Rwpos75_13 in75 sp13 11140.846016
Rwpos75_14 in75 sp14 3183.098862
Rwpos75_15 in75 sp15 3183.098862
Rwpos75_16 in75 sp16 11140.846016
Rwpos75_17 in75 sp17 3183.098862
Rwpos75_18 in75 sp18 11140.846016
Rwpos75_19 in75 sp19 3183.098862
Rwpos75_20 in75 sp20 3183.098862
Rwpos75_21 in75 sp21 11140.846016
Rwpos75_22 in75 sp22 3183.098862
Rwpos75_23 in75 sp23 3183.098862
Rwpos75_24 in75 sp24 3183.098862
Rwpos75_25 in75 sp25 11140.846016
Rwpos75_26 in75 sp26 11140.846016
Rwpos75_27 in75 sp27 3183.098862
Rwpos75_28 in75 sp28 11140.846016
Rwpos75_29 in75 sp29 11140.846016
Rwpos75_30 in75 sp30 3183.098862
Rwpos75_31 in75 sp31 3183.098862
Rwpos75_32 in75 sp32 11140.846016
Rwpos75_33 in75 sp33 3183.098862
Rwpos75_34 in75 sp34 3183.098862
Rwpos75_35 in75 sp35 11140.846016
Rwpos75_36 in75 sp36 3183.098862
Rwpos75_37 in75 sp37 3183.098862
Rwpos75_38 in75 sp38 3183.098862
Rwpos75_39 in75 sp39 3183.098862
Rwpos75_40 in75 sp40 11140.846016
Rwpos75_41 in75 sp41 11140.846016
Rwpos75_42 in75 sp42 3183.098862
Rwpos75_43 in75 sp43 3183.098862
Rwpos75_44 in75 sp44 11140.846016
Rwpos75_45 in75 sp45 3183.098862
Rwpos75_46 in75 sp46 3183.098862
Rwpos75_47 in75 sp47 11140.846016
Rwpos75_48 in75 sp48 11140.846016
Rwpos75_49 in75 sp49 3183.098862
Rwpos75_50 in75 sp50 3183.098862
Rwpos75_51 in75 sp51 3183.098862
Rwpos75_52 in75 sp52 3183.098862
Rwpos75_53 in75 sp53 3183.098862
Rwpos75_54 in75 sp54 3183.098862
Rwpos75_55 in75 sp55 3183.098862
Rwpos75_56 in75 sp56 3183.098862
Rwpos75_57 in75 sp57 11140.846016
Rwpos75_58 in75 sp58 11140.846016
Rwpos75_59 in75 sp59 3183.098862
Rwpos75_60 in75 sp60 3183.098862
Rwpos75_61 in75 sp61 11140.846016
Rwpos75_62 in75 sp62 11140.846016
Rwpos75_63 in75 sp63 3183.098862
Rwpos75_64 in75 sp64 11140.846016
Rwpos75_65 in75 sp65 3183.098862
Rwpos75_66 in75 sp66 11140.846016
Rwpos75_67 in75 sp67 11140.846016
Rwpos75_68 in75 sp68 3183.098862
Rwpos75_69 in75 sp69 3183.098862
Rwpos75_70 in75 sp70 3183.098862
Rwpos75_71 in75 sp71 11140.846016
Rwpos75_72 in75 sp72 3183.098862
Rwpos75_73 in75 sp73 11140.846016
Rwpos75_74 in75 sp74 3183.098862
Rwpos75_75 in75 sp75 3183.098862
Rwpos75_76 in75 sp76 11140.846016
Rwpos75_77 in75 sp77 3183.098862
Rwpos75_78 in75 sp78 11140.846016
Rwpos75_79 in75 sp79 3183.098862
Rwpos75_80 in75 sp80 3183.098862
Rwpos75_81 in75 sp81 11140.846016
Rwpos75_82 in75 sp82 11140.846016
Rwpos75_83 in75 sp83 3183.098862
Rwpos75_84 in75 sp84 3183.098862
Rwpos75_85 in75 sp85 3183.098862
Rwpos75_86 in75 sp86 3183.098862
Rwpos75_87 in75 sp87 11140.846016
Rwpos75_88 in75 sp88 3183.098862
Rwpos75_89 in75 sp89 11140.846016
Rwpos75_90 in75 sp90 11140.846016
Rwpos75_91 in75 sp91 3183.098862
Rwpos75_92 in75 sp92 3183.098862
Rwpos75_93 in75 sp93 3183.098862
Rwpos75_94 in75 sp94 11140.846016
Rwpos75_95 in75 sp95 3183.098862
Rwpos75_96 in75 sp96 11140.846016
Rwpos75_97 in75 sp97 11140.846016
Rwpos75_98 in75 sp98 11140.846016
Rwpos75_99 in75 sp99 3183.098862
Rwpos75_100 in75 sp100 11140.846016
Rwpos76_1 in76 sp1 3183.098862
Rwpos76_2 in76 sp2 3183.098862
Rwpos76_3 in76 sp3 11140.846016
Rwpos76_4 in76 sp4 11140.846016
Rwpos76_5 in76 sp5 11140.846016
Rwpos76_6 in76 sp6 3183.098862
Rwpos76_7 in76 sp7 3183.098862
Rwpos76_8 in76 sp8 11140.846016
Rwpos76_9 in76 sp9 3183.098862
Rwpos76_10 in76 sp10 11140.846016
Rwpos76_11 in76 sp11 3183.098862
Rwpos76_12 in76 sp12 11140.846016
Rwpos76_13 in76 sp13 3183.098862
Rwpos76_14 in76 sp14 3183.098862
Rwpos76_15 in76 sp15 11140.846016
Rwpos76_16 in76 sp16 11140.846016
Rwpos76_17 in76 sp17 3183.098862
Rwpos76_18 in76 sp18 3183.098862
Rwpos76_19 in76 sp19 11140.846016
Rwpos76_20 in76 sp20 11140.846016
Rwpos76_21 in76 sp21 11140.846016
Rwpos76_22 in76 sp22 11140.846016
Rwpos76_23 in76 sp23 3183.098862
Rwpos76_24 in76 sp24 3183.098862
Rwpos76_25 in76 sp25 3183.098862
Rwpos76_26 in76 sp26 11140.846016
Rwpos76_27 in76 sp27 11140.846016
Rwpos76_28 in76 sp28 3183.098862
Rwpos76_29 in76 sp29 11140.846016
Rwpos76_30 in76 sp30 11140.846016
Rwpos76_31 in76 sp31 3183.098862
Rwpos76_32 in76 sp32 3183.098862
Rwpos76_33 in76 sp33 3183.098862
Rwpos76_34 in76 sp34 3183.098862
Rwpos76_35 in76 sp35 11140.846016
Rwpos76_36 in76 sp36 11140.846016
Rwpos76_37 in76 sp37 3183.098862
Rwpos76_38 in76 sp38 3183.098862
Rwpos76_39 in76 sp39 3183.098862
Rwpos76_40 in76 sp40 3183.098862
Rwpos76_41 in76 sp41 11140.846016
Rwpos76_42 in76 sp42 11140.846016
Rwpos76_43 in76 sp43 3183.098862
Rwpos76_44 in76 sp44 11140.846016
Rwpos76_45 in76 sp45 11140.846016
Rwpos76_46 in76 sp46 3183.098862
Rwpos76_47 in76 sp47 3183.098862
Rwpos76_48 in76 sp48 11140.846016
Rwpos76_49 in76 sp49 3183.098862
Rwpos76_50 in76 sp50 3183.098862
Rwpos76_51 in76 sp51 11140.846016
Rwpos76_52 in76 sp52 3183.098862
Rwpos76_53 in76 sp53 3183.098862
Rwpos76_54 in76 sp54 11140.846016
Rwpos76_55 in76 sp55 11140.846016
Rwpos76_56 in76 sp56 11140.846016
Rwpos76_57 in76 sp57 3183.098862
Rwpos76_58 in76 sp58 11140.846016
Rwpos76_59 in76 sp59 3183.098862
Rwpos76_60 in76 sp60 11140.846016
Rwpos76_61 in76 sp61 11140.846016
Rwpos76_62 in76 sp62 3183.098862
Rwpos76_63 in76 sp63 11140.846016
Rwpos76_64 in76 sp64 11140.846016
Rwpos76_65 in76 sp65 3183.098862
Rwpos76_66 in76 sp66 11140.846016
Rwpos76_67 in76 sp67 3183.098862
Rwpos76_68 in76 sp68 11140.846016
Rwpos76_69 in76 sp69 3183.098862
Rwpos76_70 in76 sp70 3183.098862
Rwpos76_71 in76 sp71 3183.098862
Rwpos76_72 in76 sp72 3183.098862
Rwpos76_73 in76 sp73 11140.846016
Rwpos76_74 in76 sp74 3183.098862
Rwpos76_75 in76 sp75 3183.098862
Rwpos76_76 in76 sp76 3183.098862
Rwpos76_77 in76 sp77 3183.098862
Rwpos76_78 in76 sp78 3183.098862
Rwpos76_79 in76 sp79 11140.846016
Rwpos76_80 in76 sp80 3183.098862
Rwpos76_81 in76 sp81 11140.846016
Rwpos76_82 in76 sp82 11140.846016
Rwpos76_83 in76 sp83 3183.098862
Rwpos76_84 in76 sp84 11140.846016
Rwpos76_85 in76 sp85 3183.098862
Rwpos76_86 in76 sp86 3183.098862
Rwpos76_87 in76 sp87 11140.846016
Rwpos76_88 in76 sp88 3183.098862
Rwpos76_89 in76 sp89 3183.098862
Rwpos76_90 in76 sp90 3183.098862
Rwpos76_91 in76 sp91 3183.098862
Rwpos76_92 in76 sp92 3183.098862
Rwpos76_93 in76 sp93 11140.846016
Rwpos76_94 in76 sp94 11140.846016
Rwpos76_95 in76 sp95 3183.098862
Rwpos76_96 in76 sp96 11140.846016
Rwpos76_97 in76 sp97 3183.098862
Rwpos76_98 in76 sp98 11140.846016
Rwpos76_99 in76 sp99 3183.098862
Rwpos76_100 in76 sp100 3183.098862
Rwpos77_1 in77 sp1 11140.846016
Rwpos77_2 in77 sp2 3183.098862
Rwpos77_3 in77 sp3 11140.846016
Rwpos77_4 in77 sp4 3183.098862
Rwpos77_5 in77 sp5 3183.098862
Rwpos77_6 in77 sp6 11140.846016
Rwpos77_7 in77 sp7 11140.846016
Rwpos77_8 in77 sp8 11140.846016
Rwpos77_9 in77 sp9 3183.098862
Rwpos77_10 in77 sp10 3183.098862
Rwpos77_11 in77 sp11 11140.846016
Rwpos77_12 in77 sp12 3183.098862
Rwpos77_13 in77 sp13 3183.098862
Rwpos77_14 in77 sp14 3183.098862
Rwpos77_15 in77 sp15 11140.846016
Rwpos77_16 in77 sp16 3183.098862
Rwpos77_17 in77 sp17 3183.098862
Rwpos77_18 in77 sp18 11140.846016
Rwpos77_19 in77 sp19 3183.098862
Rwpos77_20 in77 sp20 11140.846016
Rwpos77_21 in77 sp21 11140.846016
Rwpos77_22 in77 sp22 11140.846016
Rwpos77_23 in77 sp23 11140.846016
Rwpos77_24 in77 sp24 11140.846016
Rwpos77_25 in77 sp25 3183.098862
Rwpos77_26 in77 sp26 11140.846016
Rwpos77_27 in77 sp27 3183.098862
Rwpos77_28 in77 sp28 11140.846016
Rwpos77_29 in77 sp29 3183.098862
Rwpos77_30 in77 sp30 11140.846016
Rwpos77_31 in77 sp31 3183.098862
Rwpos77_32 in77 sp32 11140.846016
Rwpos77_33 in77 sp33 11140.846016
Rwpos77_34 in77 sp34 3183.098862
Rwpos77_35 in77 sp35 3183.098862
Rwpos77_36 in77 sp36 11140.846016
Rwpos77_37 in77 sp37 11140.846016
Rwpos77_38 in77 sp38 11140.846016
Rwpos77_39 in77 sp39 3183.098862
Rwpos77_40 in77 sp40 3183.098862
Rwpos77_41 in77 sp41 11140.846016
Rwpos77_42 in77 sp42 3183.098862
Rwpos77_43 in77 sp43 11140.846016
Rwpos77_44 in77 sp44 11140.846016
Rwpos77_45 in77 sp45 11140.846016
Rwpos77_46 in77 sp46 3183.098862
Rwpos77_47 in77 sp47 11140.846016
Rwpos77_48 in77 sp48 3183.098862
Rwpos77_49 in77 sp49 3183.098862
Rwpos77_50 in77 sp50 3183.098862
Rwpos77_51 in77 sp51 3183.098862
Rwpos77_52 in77 sp52 3183.098862
Rwpos77_53 in77 sp53 11140.846016
Rwpos77_54 in77 sp54 3183.098862
Rwpos77_55 in77 sp55 3183.098862
Rwpos77_56 in77 sp56 3183.098862
Rwpos77_57 in77 sp57 3183.098862
Rwpos77_58 in77 sp58 3183.098862
Rwpos77_59 in77 sp59 11140.846016
Rwpos77_60 in77 sp60 3183.098862
Rwpos77_61 in77 sp61 11140.846016
Rwpos77_62 in77 sp62 3183.098862
Rwpos77_63 in77 sp63 3183.098862
Rwpos77_64 in77 sp64 11140.846016
Rwpos77_65 in77 sp65 3183.098862
Rwpos77_66 in77 sp66 3183.098862
Rwpos77_67 in77 sp67 11140.846016
Rwpos77_68 in77 sp68 11140.846016
Rwpos77_69 in77 sp69 3183.098862
Rwpos77_70 in77 sp70 11140.846016
Rwpos77_71 in77 sp71 3183.098862
Rwpos77_72 in77 sp72 3183.098862
Rwpos77_73 in77 sp73 3183.098862
Rwpos77_74 in77 sp74 11140.846016
Rwpos77_75 in77 sp75 11140.846016
Rwpos77_76 in77 sp76 11140.846016
Rwpos77_77 in77 sp77 3183.098862
Rwpos77_78 in77 sp78 3183.098862
Rwpos77_79 in77 sp79 3183.098862
Rwpos77_80 in77 sp80 3183.098862
Rwpos77_81 in77 sp81 11140.846016
Rwpos77_82 in77 sp82 3183.098862
Rwpos77_83 in77 sp83 3183.098862
Rwpos77_84 in77 sp84 3183.098862
Rwpos77_85 in77 sp85 3183.098862
Rwpos77_86 in77 sp86 3183.098862
Rwpos77_87 in77 sp87 3183.098862
Rwpos77_88 in77 sp88 3183.098862
Rwpos77_89 in77 sp89 11140.846016
Rwpos77_90 in77 sp90 11140.846016
Rwpos77_91 in77 sp91 11140.846016
Rwpos77_92 in77 sp92 11140.846016
Rwpos77_93 in77 sp93 3183.098862
Rwpos77_94 in77 sp94 11140.846016
Rwpos77_95 in77 sp95 3183.098862
Rwpos77_96 in77 sp96 11140.846016
Rwpos77_97 in77 sp97 11140.846016
Rwpos77_98 in77 sp98 3183.098862
Rwpos77_99 in77 sp99 3183.098862
Rwpos77_100 in77 sp100 11140.846016
Rwpos78_1 in78 sp1 3183.098862
Rwpos78_2 in78 sp2 3183.098862
Rwpos78_3 in78 sp3 3183.098862
Rwpos78_4 in78 sp4 3183.098862
Rwpos78_5 in78 sp5 11140.846016
Rwpos78_6 in78 sp6 3183.098862
Rwpos78_7 in78 sp7 11140.846016
Rwpos78_8 in78 sp8 11140.846016
Rwpos78_9 in78 sp9 3183.098862
Rwpos78_10 in78 sp10 3183.098862
Rwpos78_11 in78 sp11 11140.846016
Rwpos78_12 in78 sp12 11140.846016
Rwpos78_13 in78 sp13 3183.098862
Rwpos78_14 in78 sp14 3183.098862
Rwpos78_15 in78 sp15 3183.098862
Rwpos78_16 in78 sp16 3183.098862
Rwpos78_17 in78 sp17 3183.098862
Rwpos78_18 in78 sp18 3183.098862
Rwpos78_19 in78 sp19 11140.846016
Rwpos78_20 in78 sp20 11140.846016
Rwpos78_21 in78 sp21 11140.846016
Rwpos78_22 in78 sp22 11140.846016
Rwpos78_23 in78 sp23 11140.846016
Rwpos78_24 in78 sp24 11140.846016
Rwpos78_25 in78 sp25 3183.098862
Rwpos78_26 in78 sp26 3183.098862
Rwpos78_27 in78 sp27 11140.846016
Rwpos78_28 in78 sp28 11140.846016
Rwpos78_29 in78 sp29 3183.098862
Rwpos78_30 in78 sp30 11140.846016
Rwpos78_31 in78 sp31 11140.846016
Rwpos78_32 in78 sp32 3183.098862
Rwpos78_33 in78 sp33 3183.098862
Rwpos78_34 in78 sp34 3183.098862
Rwpos78_35 in78 sp35 11140.846016
Rwpos78_36 in78 sp36 11140.846016
Rwpos78_37 in78 sp37 3183.098862
Rwpos78_38 in78 sp38 11140.846016
Rwpos78_39 in78 sp39 11140.846016
Rwpos78_40 in78 sp40 11140.846016
Rwpos78_41 in78 sp41 3183.098862
Rwpos78_42 in78 sp42 3183.098862
Rwpos78_43 in78 sp43 11140.846016
Rwpos78_44 in78 sp44 3183.098862
Rwpos78_45 in78 sp45 3183.098862
Rwpos78_46 in78 sp46 3183.098862
Rwpos78_47 in78 sp47 11140.846016
Rwpos78_48 in78 sp48 3183.098862
Rwpos78_49 in78 sp49 11140.846016
Rwpos78_50 in78 sp50 3183.098862
Rwpos78_51 in78 sp51 3183.098862
Rwpos78_52 in78 sp52 11140.846016
Rwpos78_53 in78 sp53 11140.846016
Rwpos78_54 in78 sp54 11140.846016
Rwpos78_55 in78 sp55 3183.098862
Rwpos78_56 in78 sp56 3183.098862
Rwpos78_57 in78 sp57 3183.098862
Rwpos78_58 in78 sp58 3183.098862
Rwpos78_59 in78 sp59 11140.846016
Rwpos78_60 in78 sp60 11140.846016
Rwpos78_61 in78 sp61 3183.098862
Rwpos78_62 in78 sp62 11140.846016
Rwpos78_63 in78 sp63 11140.846016
Rwpos78_64 in78 sp64 3183.098862
Rwpos78_65 in78 sp65 3183.098862
Rwpos78_66 in78 sp66 3183.098862
Rwpos78_67 in78 sp67 3183.098862
Rwpos78_68 in78 sp68 11140.846016
Rwpos78_69 in78 sp69 3183.098862
Rwpos78_70 in78 sp70 11140.846016
Rwpos78_71 in78 sp71 3183.098862
Rwpos78_72 in78 sp72 3183.098862
Rwpos78_73 in78 sp73 3183.098862
Rwpos78_74 in78 sp74 11140.846016
Rwpos78_75 in78 sp75 11140.846016
Rwpos78_76 in78 sp76 11140.846016
Rwpos78_77 in78 sp77 3183.098862
Rwpos78_78 in78 sp78 11140.846016
Rwpos78_79 in78 sp79 11140.846016
Rwpos78_80 in78 sp80 3183.098862
Rwpos78_81 in78 sp81 3183.098862
Rwpos78_82 in78 sp82 3183.098862
Rwpos78_83 in78 sp83 3183.098862
Rwpos78_84 in78 sp84 3183.098862
Rwpos78_85 in78 sp85 3183.098862
Rwpos78_86 in78 sp86 3183.098862
Rwpos78_87 in78 sp87 3183.098862
Rwpos78_88 in78 sp88 11140.846016
Rwpos78_89 in78 sp89 3183.098862
Rwpos78_90 in78 sp90 11140.846016
Rwpos78_91 in78 sp91 3183.098862
Rwpos78_92 in78 sp92 11140.846016
Rwpos78_93 in78 sp93 3183.098862
Rwpos78_94 in78 sp94 11140.846016
Rwpos78_95 in78 sp95 11140.846016
Rwpos78_96 in78 sp96 3183.098862
Rwpos78_97 in78 sp97 3183.098862
Rwpos78_98 in78 sp98 3183.098862
Rwpos78_99 in78 sp99 3183.098862
Rwpos78_100 in78 sp100 11140.846016
Rwpos79_1 in79 sp1 3183.098862
Rwpos79_2 in79 sp2 11140.846016
Rwpos79_3 in79 sp3 3183.098862
Rwpos79_4 in79 sp4 11140.846016
Rwpos79_5 in79 sp5 11140.846016
Rwpos79_6 in79 sp6 11140.846016
Rwpos79_7 in79 sp7 3183.098862
Rwpos79_8 in79 sp8 11140.846016
Rwpos79_9 in79 sp9 3183.098862
Rwpos79_10 in79 sp10 11140.846016
Rwpos79_11 in79 sp11 11140.846016
Rwpos79_12 in79 sp12 11140.846016
Rwpos79_13 in79 sp13 11140.846016
Rwpos79_14 in79 sp14 3183.098862
Rwpos79_15 in79 sp15 3183.098862
Rwpos79_16 in79 sp16 3183.098862
Rwpos79_17 in79 sp17 3183.098862
Rwpos79_18 in79 sp18 11140.846016
Rwpos79_19 in79 sp19 3183.098862
Rwpos79_20 in79 sp20 3183.098862
Rwpos79_21 in79 sp21 11140.846016
Rwpos79_22 in79 sp22 11140.846016
Rwpos79_23 in79 sp23 3183.098862
Rwpos79_24 in79 sp24 11140.846016
Rwpos79_25 in79 sp25 3183.098862
Rwpos79_26 in79 sp26 11140.846016
Rwpos79_27 in79 sp27 3183.098862
Rwpos79_28 in79 sp28 11140.846016
Rwpos79_29 in79 sp29 11140.846016
Rwpos79_30 in79 sp30 3183.098862
Rwpos79_31 in79 sp31 11140.846016
Rwpos79_32 in79 sp32 11140.846016
Rwpos79_33 in79 sp33 3183.098862
Rwpos79_34 in79 sp34 11140.846016
Rwpos79_35 in79 sp35 11140.846016
Rwpos79_36 in79 sp36 3183.098862
Rwpos79_37 in79 sp37 11140.846016
Rwpos79_38 in79 sp38 11140.846016
Rwpos79_39 in79 sp39 3183.098862
Rwpos79_40 in79 sp40 11140.846016
Rwpos79_41 in79 sp41 3183.098862
Rwpos79_42 in79 sp42 11140.846016
Rwpos79_43 in79 sp43 3183.098862
Rwpos79_44 in79 sp44 11140.846016
Rwpos79_45 in79 sp45 11140.846016
Rwpos79_46 in79 sp46 3183.098862
Rwpos79_47 in79 sp47 11140.846016
Rwpos79_48 in79 sp48 11140.846016
Rwpos79_49 in79 sp49 3183.098862
Rwpos79_50 in79 sp50 11140.846016
Rwpos79_51 in79 sp51 11140.846016
Rwpos79_52 in79 sp52 3183.098862
Rwpos79_53 in79 sp53 3183.098862
Rwpos79_54 in79 sp54 11140.846016
Rwpos79_55 in79 sp55 3183.098862
Rwpos79_56 in79 sp56 11140.846016
Rwpos79_57 in79 sp57 3183.098862
Rwpos79_58 in79 sp58 3183.098862
Rwpos79_59 in79 sp59 3183.098862
Rwpos79_60 in79 sp60 11140.846016
Rwpos79_61 in79 sp61 11140.846016
Rwpos79_62 in79 sp62 3183.098862
Rwpos79_63 in79 sp63 3183.098862
Rwpos79_64 in79 sp64 11140.846016
Rwpos79_65 in79 sp65 3183.098862
Rwpos79_66 in79 sp66 11140.846016
Rwpos79_67 in79 sp67 11140.846016
Rwpos79_68 in79 sp68 11140.846016
Rwpos79_69 in79 sp69 3183.098862
Rwpos79_70 in79 sp70 3183.098862
Rwpos79_71 in79 sp71 3183.098862
Rwpos79_72 in79 sp72 11140.846016
Rwpos79_73 in79 sp73 11140.846016
Rwpos79_74 in79 sp74 3183.098862
Rwpos79_75 in79 sp75 11140.846016
Rwpos79_76 in79 sp76 3183.098862
Rwpos79_77 in79 sp77 11140.846016
Rwpos79_78 in79 sp78 3183.098862
Rwpos79_79 in79 sp79 3183.098862
Rwpos79_80 in79 sp80 11140.846016
Rwpos79_81 in79 sp81 3183.098862
Rwpos79_82 in79 sp82 11140.846016
Rwpos79_83 in79 sp83 11140.846016
Rwpos79_84 in79 sp84 3183.098862
Rwpos79_85 in79 sp85 11140.846016
Rwpos79_86 in79 sp86 3183.098862
Rwpos79_87 in79 sp87 3183.098862
Rwpos79_88 in79 sp88 3183.098862
Rwpos79_89 in79 sp89 11140.846016
Rwpos79_90 in79 sp90 11140.846016
Rwpos79_91 in79 sp91 11140.846016
Rwpos79_92 in79 sp92 11140.846016
Rwpos79_93 in79 sp93 11140.846016
Rwpos79_94 in79 sp94 3183.098862
Rwpos79_95 in79 sp95 3183.098862
Rwpos79_96 in79 sp96 11140.846016
Rwpos79_97 in79 sp97 3183.098862
Rwpos79_98 in79 sp98 3183.098862
Rwpos79_99 in79 sp99 11140.846016
Rwpos79_100 in79 sp100 11140.846016
Rwpos80_1 in80 sp1 3183.098862
Rwpos80_2 in80 sp2 3183.098862
Rwpos80_3 in80 sp3 11140.846016
Rwpos80_4 in80 sp4 11140.846016
Rwpos80_5 in80 sp5 11140.846016
Rwpos80_6 in80 sp6 3183.098862
Rwpos80_7 in80 sp7 3183.098862
Rwpos80_8 in80 sp8 3183.098862
Rwpos80_9 in80 sp9 11140.846016
Rwpos80_10 in80 sp10 11140.846016
Rwpos80_11 in80 sp11 11140.846016
Rwpos80_12 in80 sp12 3183.098862
Rwpos80_13 in80 sp13 11140.846016
Rwpos80_14 in80 sp14 11140.846016
Rwpos80_15 in80 sp15 11140.846016
Rwpos80_16 in80 sp16 11140.846016
Rwpos80_17 in80 sp17 11140.846016
Rwpos80_18 in80 sp18 3183.098862
Rwpos80_19 in80 sp19 3183.098862
Rwpos80_20 in80 sp20 3183.098862
Rwpos80_21 in80 sp21 11140.846016
Rwpos80_22 in80 sp22 3183.098862
Rwpos80_23 in80 sp23 3183.098862
Rwpos80_24 in80 sp24 3183.098862
Rwpos80_25 in80 sp25 11140.846016
Rwpos80_26 in80 sp26 11140.846016
Rwpos80_27 in80 sp27 3183.098862
Rwpos80_28 in80 sp28 11140.846016
Rwpos80_29 in80 sp29 11140.846016
Rwpos80_30 in80 sp30 3183.098862
Rwpos80_31 in80 sp31 11140.846016
Rwpos80_32 in80 sp32 3183.098862
Rwpos80_33 in80 sp33 11140.846016
Rwpos80_34 in80 sp34 3183.098862
Rwpos80_35 in80 sp35 11140.846016
Rwpos80_36 in80 sp36 11140.846016
Rwpos80_37 in80 sp37 11140.846016
Rwpos80_38 in80 sp38 3183.098862
Rwpos80_39 in80 sp39 3183.098862
Rwpos80_40 in80 sp40 11140.846016
Rwpos80_41 in80 sp41 3183.098862
Rwpos80_42 in80 sp42 11140.846016
Rwpos80_43 in80 sp43 3183.098862
Rwpos80_44 in80 sp44 3183.098862
Rwpos80_45 in80 sp45 3183.098862
Rwpos80_46 in80 sp46 11140.846016
Rwpos80_47 in80 sp47 11140.846016
Rwpos80_48 in80 sp48 3183.098862
Rwpos80_49 in80 sp49 3183.098862
Rwpos80_50 in80 sp50 3183.098862
Rwpos80_51 in80 sp51 3183.098862
Rwpos80_52 in80 sp52 11140.846016
Rwpos80_53 in80 sp53 11140.846016
Rwpos80_54 in80 sp54 3183.098862
Rwpos80_55 in80 sp55 3183.098862
Rwpos80_56 in80 sp56 3183.098862
Rwpos80_57 in80 sp57 11140.846016
Rwpos80_58 in80 sp58 11140.846016
Rwpos80_59 in80 sp59 3183.098862
Rwpos80_60 in80 sp60 3183.098862
Rwpos80_61 in80 sp61 11140.846016
Rwpos80_62 in80 sp62 11140.846016
Rwpos80_63 in80 sp63 11140.846016
Rwpos80_64 in80 sp64 3183.098862
Rwpos80_65 in80 sp65 3183.098862
Rwpos80_66 in80 sp66 3183.098862
Rwpos80_67 in80 sp67 3183.098862
Rwpos80_68 in80 sp68 11140.846016
Rwpos80_69 in80 sp69 11140.846016
Rwpos80_70 in80 sp70 3183.098862
Rwpos80_71 in80 sp71 3183.098862
Rwpos80_72 in80 sp72 3183.098862
Rwpos80_73 in80 sp73 11140.846016
Rwpos80_74 in80 sp74 11140.846016
Rwpos80_75 in80 sp75 3183.098862
Rwpos80_76 in80 sp76 3183.098862
Rwpos80_77 in80 sp77 11140.846016
Rwpos80_78 in80 sp78 11140.846016
Rwpos80_79 in80 sp79 11140.846016
Rwpos80_80 in80 sp80 11140.846016
Rwpos80_81 in80 sp81 3183.098862
Rwpos80_82 in80 sp82 3183.098862
Rwpos80_83 in80 sp83 11140.846016
Rwpos80_84 in80 sp84 3183.098862
Rwpos80_85 in80 sp85 3183.098862
Rwpos80_86 in80 sp86 3183.098862
Rwpos80_87 in80 sp87 3183.098862
Rwpos80_88 in80 sp88 3183.098862
Rwpos80_89 in80 sp89 3183.098862
Rwpos80_90 in80 sp90 3183.098862
Rwpos80_91 in80 sp91 11140.846016
Rwpos80_92 in80 sp92 3183.098862
Rwpos80_93 in80 sp93 3183.098862
Rwpos80_94 in80 sp94 11140.846016
Rwpos80_95 in80 sp95 3183.098862
Rwpos80_96 in80 sp96 3183.098862
Rwpos80_97 in80 sp97 3183.098862
Rwpos80_98 in80 sp98 3183.098862
Rwpos80_99 in80 sp99 11140.846016
Rwpos80_100 in80 sp100 11140.846016
Rwpos81_1 in81 sp1 3183.098862
Rwpos81_2 in81 sp2 11140.846016
Rwpos81_3 in81 sp3 11140.846016
Rwpos81_4 in81 sp4 3183.098862
Rwpos81_5 in81 sp5 11140.846016
Rwpos81_6 in81 sp6 11140.846016
Rwpos81_7 in81 sp7 3183.098862
Rwpos81_8 in81 sp8 3183.098862
Rwpos81_9 in81 sp9 11140.846016
Rwpos81_10 in81 sp10 3183.098862
Rwpos81_11 in81 sp11 11140.846016
Rwpos81_12 in81 sp12 3183.098862
Rwpos81_13 in81 sp13 11140.846016
Rwpos81_14 in81 sp14 11140.846016
Rwpos81_15 in81 sp15 11140.846016
Rwpos81_16 in81 sp16 3183.098862
Rwpos81_17 in81 sp17 3183.098862
Rwpos81_18 in81 sp18 3183.098862
Rwpos81_19 in81 sp19 3183.098862
Rwpos81_20 in81 sp20 3183.098862
Rwpos81_21 in81 sp21 11140.846016
Rwpos81_22 in81 sp22 3183.098862
Rwpos81_23 in81 sp23 11140.846016
Rwpos81_24 in81 sp24 3183.098862
Rwpos81_25 in81 sp25 3183.098862
Rwpos81_26 in81 sp26 3183.098862
Rwpos81_27 in81 sp27 11140.846016
Rwpos81_28 in81 sp28 3183.098862
Rwpos81_29 in81 sp29 3183.098862
Rwpos81_30 in81 sp30 3183.098862
Rwpos81_31 in81 sp31 11140.846016
Rwpos81_32 in81 sp32 11140.846016
Rwpos81_33 in81 sp33 11140.846016
Rwpos81_34 in81 sp34 11140.846016
Rwpos81_35 in81 sp35 11140.846016
Rwpos81_36 in81 sp36 3183.098862
Rwpos81_37 in81 sp37 11140.846016
Rwpos81_38 in81 sp38 11140.846016
Rwpos81_39 in81 sp39 11140.846016
Rwpos81_40 in81 sp40 3183.098862
Rwpos81_41 in81 sp41 3183.098862
Rwpos81_42 in81 sp42 3183.098862
Rwpos81_43 in81 sp43 3183.098862
Rwpos81_44 in81 sp44 11140.846016
Rwpos81_45 in81 sp45 3183.098862
Rwpos81_46 in81 sp46 11140.846016
Rwpos81_47 in81 sp47 11140.846016
Rwpos81_48 in81 sp48 11140.846016
Rwpos81_49 in81 sp49 3183.098862
Rwpos81_50 in81 sp50 11140.846016
Rwpos81_51 in81 sp51 3183.098862
Rwpos81_52 in81 sp52 3183.098862
Rwpos81_53 in81 sp53 11140.846016
Rwpos81_54 in81 sp54 3183.098862
Rwpos81_55 in81 sp55 11140.846016
Rwpos81_56 in81 sp56 11140.846016
Rwpos81_57 in81 sp57 11140.846016
Rwpos81_58 in81 sp58 11140.846016
Rwpos81_59 in81 sp59 3183.098862
Rwpos81_60 in81 sp60 11140.846016
Rwpos81_61 in81 sp61 11140.846016
Rwpos81_62 in81 sp62 11140.846016
Rwpos81_63 in81 sp63 3183.098862
Rwpos81_64 in81 sp64 11140.846016
Rwpos81_65 in81 sp65 3183.098862
Rwpos81_66 in81 sp66 3183.098862
Rwpos81_67 in81 sp67 3183.098862
Rwpos81_68 in81 sp68 3183.098862
Rwpos81_69 in81 sp69 3183.098862
Rwpos81_70 in81 sp70 3183.098862
Rwpos81_71 in81 sp71 11140.846016
Rwpos81_72 in81 sp72 3183.098862
Rwpos81_73 in81 sp73 3183.098862
Rwpos81_74 in81 sp74 11140.846016
Rwpos81_75 in81 sp75 3183.098862
Rwpos81_76 in81 sp76 3183.098862
Rwpos81_77 in81 sp77 11140.846016
Rwpos81_78 in81 sp78 11140.846016
Rwpos81_79 in81 sp79 11140.846016
Rwpos81_80 in81 sp80 11140.846016
Rwpos81_81 in81 sp81 3183.098862
Rwpos81_82 in81 sp82 11140.846016
Rwpos81_83 in81 sp83 3183.098862
Rwpos81_84 in81 sp84 3183.098862
Rwpos81_85 in81 sp85 3183.098862
Rwpos81_86 in81 sp86 3183.098862
Rwpos81_87 in81 sp87 3183.098862
Rwpos81_88 in81 sp88 11140.846016
Rwpos81_89 in81 sp89 11140.846016
Rwpos81_90 in81 sp90 3183.098862
Rwpos81_91 in81 sp91 3183.098862
Rwpos81_92 in81 sp92 11140.846016
Rwpos81_93 in81 sp93 11140.846016
Rwpos81_94 in81 sp94 11140.846016
Rwpos81_95 in81 sp95 3183.098862
Rwpos81_96 in81 sp96 11140.846016
Rwpos81_97 in81 sp97 11140.846016
Rwpos81_98 in81 sp98 11140.846016
Rwpos81_99 in81 sp99 11140.846016
Rwpos81_100 in81 sp100 11140.846016
Rwpos82_1 in82 sp1 11140.846016
Rwpos82_2 in82 sp2 3183.098862
Rwpos82_3 in82 sp3 11140.846016
Rwpos82_4 in82 sp4 3183.098862
Rwpos82_5 in82 sp5 11140.846016
Rwpos82_6 in82 sp6 11140.846016
Rwpos82_7 in82 sp7 3183.098862
Rwpos82_8 in82 sp8 3183.098862
Rwpos82_9 in82 sp9 3183.098862
Rwpos82_10 in82 sp10 3183.098862
Rwpos82_11 in82 sp11 11140.846016
Rwpos82_12 in82 sp12 11140.846016
Rwpos82_13 in82 sp13 11140.846016
Rwpos82_14 in82 sp14 3183.098862
Rwpos82_15 in82 sp15 11140.846016
Rwpos82_16 in82 sp16 3183.098862
Rwpos82_17 in82 sp17 11140.846016
Rwpos82_18 in82 sp18 11140.846016
Rwpos82_19 in82 sp19 3183.098862
Rwpos82_20 in82 sp20 11140.846016
Rwpos82_21 in82 sp21 11140.846016
Rwpos82_22 in82 sp22 11140.846016
Rwpos82_23 in82 sp23 3183.098862
Rwpos82_24 in82 sp24 3183.098862
Rwpos82_25 in82 sp25 3183.098862
Rwpos82_26 in82 sp26 3183.098862
Rwpos82_27 in82 sp27 3183.098862
Rwpos82_28 in82 sp28 11140.846016
Rwpos82_29 in82 sp29 11140.846016
Rwpos82_30 in82 sp30 3183.098862
Rwpos82_31 in82 sp31 11140.846016
Rwpos82_32 in82 sp32 11140.846016
Rwpos82_33 in82 sp33 11140.846016
Rwpos82_34 in82 sp34 11140.846016
Rwpos82_35 in82 sp35 3183.098862
Rwpos82_36 in82 sp36 11140.846016
Rwpos82_37 in82 sp37 3183.098862
Rwpos82_38 in82 sp38 3183.098862
Rwpos82_39 in82 sp39 11140.846016
Rwpos82_40 in82 sp40 11140.846016
Rwpos82_41 in82 sp41 11140.846016
Rwpos82_42 in82 sp42 11140.846016
Rwpos82_43 in82 sp43 11140.846016
Rwpos82_44 in82 sp44 3183.098862
Rwpos82_45 in82 sp45 3183.098862
Rwpos82_46 in82 sp46 11140.846016
Rwpos82_47 in82 sp47 3183.098862
Rwpos82_48 in82 sp48 3183.098862
Rwpos82_49 in82 sp49 3183.098862
Rwpos82_50 in82 sp50 3183.098862
Rwpos82_51 in82 sp51 3183.098862
Rwpos82_52 in82 sp52 11140.846016
Rwpos82_53 in82 sp53 3183.098862
Rwpos82_54 in82 sp54 3183.098862
Rwpos82_55 in82 sp55 11140.846016
Rwpos82_56 in82 sp56 11140.846016
Rwpos82_57 in82 sp57 3183.098862
Rwpos82_58 in82 sp58 3183.098862
Rwpos82_59 in82 sp59 11140.846016
Rwpos82_60 in82 sp60 11140.846016
Rwpos82_61 in82 sp61 3183.098862
Rwpos82_62 in82 sp62 3183.098862
Rwpos82_63 in82 sp63 3183.098862
Rwpos82_64 in82 sp64 3183.098862
Rwpos82_65 in82 sp65 3183.098862
Rwpos82_66 in82 sp66 11140.846016
Rwpos82_67 in82 sp67 11140.846016
Rwpos82_68 in82 sp68 3183.098862
Rwpos82_69 in82 sp69 11140.846016
Rwpos82_70 in82 sp70 3183.098862
Rwpos82_71 in82 sp71 11140.846016
Rwpos82_72 in82 sp72 11140.846016
Rwpos82_73 in82 sp73 11140.846016
Rwpos82_74 in82 sp74 3183.098862
Rwpos82_75 in82 sp75 11140.846016
Rwpos82_76 in82 sp76 11140.846016
Rwpos82_77 in82 sp77 3183.098862
Rwpos82_78 in82 sp78 11140.846016
Rwpos82_79 in82 sp79 3183.098862
Rwpos82_80 in82 sp80 3183.098862
Rwpos82_81 in82 sp81 3183.098862
Rwpos82_82 in82 sp82 11140.846016
Rwpos82_83 in82 sp83 3183.098862
Rwpos82_84 in82 sp84 3183.098862
Rwpos82_85 in82 sp85 11140.846016
Rwpos82_86 in82 sp86 3183.098862
Rwpos82_87 in82 sp87 3183.098862
Rwpos82_88 in82 sp88 11140.846016
Rwpos82_89 in82 sp89 3183.098862
Rwpos82_90 in82 sp90 11140.846016
Rwpos82_91 in82 sp91 11140.846016
Rwpos82_92 in82 sp92 11140.846016
Rwpos82_93 in82 sp93 3183.098862
Rwpos82_94 in82 sp94 11140.846016
Rwpos82_95 in82 sp95 3183.098862
Rwpos82_96 in82 sp96 3183.098862
Rwpos82_97 in82 sp97 3183.098862
Rwpos82_98 in82 sp98 3183.098862
Rwpos82_99 in82 sp99 3183.098862
Rwpos82_100 in82 sp100 3183.098862
Rwpos83_1 in83 sp1 3183.098862
Rwpos83_2 in83 sp2 11140.846016
Rwpos83_3 in83 sp3 11140.846016
Rwpos83_4 in83 sp4 11140.846016
Rwpos83_5 in83 sp5 3183.098862
Rwpos83_6 in83 sp6 11140.846016
Rwpos83_7 in83 sp7 11140.846016
Rwpos83_8 in83 sp8 11140.846016
Rwpos83_9 in83 sp9 3183.098862
Rwpos83_10 in83 sp10 11140.846016
Rwpos83_11 in83 sp11 11140.846016
Rwpos83_12 in83 sp12 11140.846016
Rwpos83_13 in83 sp13 11140.846016
Rwpos83_14 in83 sp14 3183.098862
Rwpos83_15 in83 sp15 3183.098862
Rwpos83_16 in83 sp16 3183.098862
Rwpos83_17 in83 sp17 3183.098862
Rwpos83_18 in83 sp18 11140.846016
Rwpos83_19 in83 sp19 3183.098862
Rwpos83_20 in83 sp20 11140.846016
Rwpos83_21 in83 sp21 11140.846016
Rwpos83_22 in83 sp22 11140.846016
Rwpos83_23 in83 sp23 11140.846016
Rwpos83_24 in83 sp24 11140.846016
Rwpos83_25 in83 sp25 3183.098862
Rwpos83_26 in83 sp26 11140.846016
Rwpos83_27 in83 sp27 11140.846016
Rwpos83_28 in83 sp28 11140.846016
Rwpos83_29 in83 sp29 3183.098862
Rwpos83_30 in83 sp30 11140.846016
Rwpos83_31 in83 sp31 3183.098862
Rwpos83_32 in83 sp32 3183.098862
Rwpos83_33 in83 sp33 3183.098862
Rwpos83_34 in83 sp34 11140.846016
Rwpos83_35 in83 sp35 3183.098862
Rwpos83_36 in83 sp36 11140.846016
Rwpos83_37 in83 sp37 3183.098862
Rwpos83_38 in83 sp38 11140.846016
Rwpos83_39 in83 sp39 11140.846016
Rwpos83_40 in83 sp40 11140.846016
Rwpos83_41 in83 sp41 3183.098862
Rwpos83_42 in83 sp42 11140.846016
Rwpos83_43 in83 sp43 3183.098862
Rwpos83_44 in83 sp44 11140.846016
Rwpos83_45 in83 sp45 3183.098862
Rwpos83_46 in83 sp46 3183.098862
Rwpos83_47 in83 sp47 3183.098862
Rwpos83_48 in83 sp48 3183.098862
Rwpos83_49 in83 sp49 3183.098862
Rwpos83_50 in83 sp50 3183.098862
Rwpos83_51 in83 sp51 3183.098862
Rwpos83_52 in83 sp52 11140.846016
Rwpos83_53 in83 sp53 3183.098862
Rwpos83_54 in83 sp54 11140.846016
Rwpos83_55 in83 sp55 3183.098862
Rwpos83_56 in83 sp56 11140.846016
Rwpos83_57 in83 sp57 3183.098862
Rwpos83_58 in83 sp58 11140.846016
Rwpos83_59 in83 sp59 11140.846016
Rwpos83_60 in83 sp60 11140.846016
Rwpos83_61 in83 sp61 11140.846016
Rwpos83_62 in83 sp62 3183.098862
Rwpos83_63 in83 sp63 11140.846016
Rwpos83_64 in83 sp64 3183.098862
Rwpos83_65 in83 sp65 3183.098862
Rwpos83_66 in83 sp66 11140.846016
Rwpos83_67 in83 sp67 3183.098862
Rwpos83_68 in83 sp68 3183.098862
Rwpos83_69 in83 sp69 3183.098862
Rwpos83_70 in83 sp70 11140.846016
Rwpos83_71 in83 sp71 3183.098862
Rwpos83_72 in83 sp72 11140.846016
Rwpos83_73 in83 sp73 3183.098862
Rwpos83_74 in83 sp74 3183.098862
Rwpos83_75 in83 sp75 3183.098862
Rwpos83_76 in83 sp76 11140.846016
Rwpos83_77 in83 sp77 3183.098862
Rwpos83_78 in83 sp78 3183.098862
Rwpos83_79 in83 sp79 11140.846016
Rwpos83_80 in83 sp80 3183.098862
Rwpos83_81 in83 sp81 3183.098862
Rwpos83_82 in83 sp82 11140.846016
Rwpos83_83 in83 sp83 3183.098862
Rwpos83_84 in83 sp84 11140.846016
Rwpos83_85 in83 sp85 3183.098862
Rwpos83_86 in83 sp86 11140.846016
Rwpos83_87 in83 sp87 3183.098862
Rwpos83_88 in83 sp88 11140.846016
Rwpos83_89 in83 sp89 3183.098862
Rwpos83_90 in83 sp90 3183.098862
Rwpos83_91 in83 sp91 11140.846016
Rwpos83_92 in83 sp92 11140.846016
Rwpos83_93 in83 sp93 3183.098862
Rwpos83_94 in83 sp94 3183.098862
Rwpos83_95 in83 sp95 3183.098862
Rwpos83_96 in83 sp96 11140.846016
Rwpos83_97 in83 sp97 3183.098862
Rwpos83_98 in83 sp98 3183.098862
Rwpos83_99 in83 sp99 3183.098862
Rwpos83_100 in83 sp100 3183.098862
Rwpos84_1 in84 sp1 3183.098862
Rwpos84_2 in84 sp2 11140.846016
Rwpos84_3 in84 sp3 11140.846016
Rwpos84_4 in84 sp4 11140.846016
Rwpos84_5 in84 sp5 3183.098862
Rwpos84_6 in84 sp6 11140.846016
Rwpos84_7 in84 sp7 3183.098862
Rwpos84_8 in84 sp8 3183.098862
Rwpos84_9 in84 sp9 3183.098862
Rwpos84_10 in84 sp10 3183.098862
Rwpos84_11 in84 sp11 3183.098862
Rwpos84_12 in84 sp12 11140.846016
Rwpos84_13 in84 sp13 3183.098862
Rwpos84_14 in84 sp14 3183.098862
Rwpos84_15 in84 sp15 11140.846016
Rwpos84_16 in84 sp16 3183.098862
Rwpos84_17 in84 sp17 3183.098862
Rwpos84_18 in84 sp18 3183.098862
Rwpos84_19 in84 sp19 3183.098862
Rwpos84_20 in84 sp20 11140.846016
Rwpos84_21 in84 sp21 3183.098862
Rwpos84_22 in84 sp22 3183.098862
Rwpos84_23 in84 sp23 3183.098862
Rwpos84_24 in84 sp24 3183.098862
Rwpos84_25 in84 sp25 3183.098862
Rwpos84_26 in84 sp26 11140.846016
Rwpos84_27 in84 sp27 11140.846016
Rwpos84_28 in84 sp28 3183.098862
Rwpos84_29 in84 sp29 11140.846016
Rwpos84_30 in84 sp30 3183.098862
Rwpos84_31 in84 sp31 11140.846016
Rwpos84_32 in84 sp32 11140.846016
Rwpos84_33 in84 sp33 3183.098862
Rwpos84_34 in84 sp34 3183.098862
Rwpos84_35 in84 sp35 3183.098862
Rwpos84_36 in84 sp36 11140.846016
Rwpos84_37 in84 sp37 3183.098862
Rwpos84_38 in84 sp38 3183.098862
Rwpos84_39 in84 sp39 3183.098862
Rwpos84_40 in84 sp40 3183.098862
Rwpos84_41 in84 sp41 3183.098862
Rwpos84_42 in84 sp42 11140.846016
Rwpos84_43 in84 sp43 11140.846016
Rwpos84_44 in84 sp44 3183.098862
Rwpos84_45 in84 sp45 11140.846016
Rwpos84_46 in84 sp46 11140.846016
Rwpos84_47 in84 sp47 11140.846016
Rwpos84_48 in84 sp48 3183.098862
Rwpos84_49 in84 sp49 11140.846016
Rwpos84_50 in84 sp50 3183.098862
Rwpos84_51 in84 sp51 3183.098862
Rwpos84_52 in84 sp52 11140.846016
Rwpos84_53 in84 sp53 11140.846016
Rwpos84_54 in84 sp54 3183.098862
Rwpos84_55 in84 sp55 11140.846016
Rwpos84_56 in84 sp56 3183.098862
Rwpos84_57 in84 sp57 11140.846016
Rwpos84_58 in84 sp58 11140.846016
Rwpos84_59 in84 sp59 11140.846016
Rwpos84_60 in84 sp60 3183.098862
Rwpos84_61 in84 sp61 11140.846016
Rwpos84_62 in84 sp62 3183.098862
Rwpos84_63 in84 sp63 3183.098862
Rwpos84_64 in84 sp64 11140.846016
Rwpos84_65 in84 sp65 3183.098862
Rwpos84_66 in84 sp66 3183.098862
Rwpos84_67 in84 sp67 3183.098862
Rwpos84_68 in84 sp68 11140.846016
Rwpos84_69 in84 sp69 3183.098862
Rwpos84_70 in84 sp70 3183.098862
Rwpos84_71 in84 sp71 3183.098862
Rwpos84_72 in84 sp72 3183.098862
Rwpos84_73 in84 sp73 11140.846016
Rwpos84_74 in84 sp74 11140.846016
Rwpos84_75 in84 sp75 3183.098862
Rwpos84_76 in84 sp76 3183.098862
Rwpos84_77 in84 sp77 3183.098862
Rwpos84_78 in84 sp78 3183.098862
Rwpos84_79 in84 sp79 11140.846016
Rwpos84_80 in84 sp80 11140.846016
Rwpos84_81 in84 sp81 3183.098862
Rwpos84_82 in84 sp82 3183.098862
Rwpos84_83 in84 sp83 3183.098862
Rwpos84_84 in84 sp84 11140.846016
Rwpos84_85 in84 sp85 3183.098862
Rwpos84_86 in84 sp86 3183.098862
Rwpos84_87 in84 sp87 3183.098862
Rwpos84_88 in84 sp88 3183.098862
Rwpos84_89 in84 sp89 3183.098862
Rwpos84_90 in84 sp90 11140.846016
Rwpos84_91 in84 sp91 3183.098862
Rwpos84_92 in84 sp92 3183.098862
Rwpos84_93 in84 sp93 11140.846016
Rwpos84_94 in84 sp94 3183.098862
Rwpos84_95 in84 sp95 3183.098862
Rwpos84_96 in84 sp96 3183.098862
Rwpos84_97 in84 sp97 11140.846016
Rwpos84_98 in84 sp98 3183.098862
Rwpos84_99 in84 sp99 3183.098862
Rwpos84_100 in84 sp100 3183.098862
Rwpos85_1 in85 sp1 11140.846016
Rwpos85_2 in85 sp2 3183.098862
Rwpos85_3 in85 sp3 3183.098862
Rwpos85_4 in85 sp4 3183.098862
Rwpos85_5 in85 sp5 3183.098862
Rwpos85_6 in85 sp6 11140.846016
Rwpos85_7 in85 sp7 3183.098862
Rwpos85_8 in85 sp8 3183.098862
Rwpos85_9 in85 sp9 3183.098862
Rwpos85_10 in85 sp10 3183.098862
Rwpos85_11 in85 sp11 11140.846016
Rwpos85_12 in85 sp12 11140.846016
Rwpos85_13 in85 sp13 3183.098862
Rwpos85_14 in85 sp14 11140.846016
Rwpos85_15 in85 sp15 3183.098862
Rwpos85_16 in85 sp16 11140.846016
Rwpos85_17 in85 sp17 3183.098862
Rwpos85_18 in85 sp18 3183.098862
Rwpos85_19 in85 sp19 11140.846016
Rwpos85_20 in85 sp20 3183.098862
Rwpos85_21 in85 sp21 3183.098862
Rwpos85_22 in85 sp22 11140.846016
Rwpos85_23 in85 sp23 11140.846016
Rwpos85_24 in85 sp24 3183.098862
Rwpos85_25 in85 sp25 11140.846016
Rwpos85_26 in85 sp26 3183.098862
Rwpos85_27 in85 sp27 11140.846016
Rwpos85_28 in85 sp28 11140.846016
Rwpos85_29 in85 sp29 11140.846016
Rwpos85_30 in85 sp30 3183.098862
Rwpos85_31 in85 sp31 3183.098862
Rwpos85_32 in85 sp32 11140.846016
Rwpos85_33 in85 sp33 3183.098862
Rwpos85_34 in85 sp34 3183.098862
Rwpos85_35 in85 sp35 11140.846016
Rwpos85_36 in85 sp36 3183.098862
Rwpos85_37 in85 sp37 3183.098862
Rwpos85_38 in85 sp38 3183.098862
Rwpos85_39 in85 sp39 3183.098862
Rwpos85_40 in85 sp40 3183.098862
Rwpos85_41 in85 sp41 11140.846016
Rwpos85_42 in85 sp42 3183.098862
Rwpos85_43 in85 sp43 11140.846016
Rwpos85_44 in85 sp44 11140.846016
Rwpos85_45 in85 sp45 11140.846016
Rwpos85_46 in85 sp46 3183.098862
Rwpos85_47 in85 sp47 3183.098862
Rwpos85_48 in85 sp48 11140.846016
Rwpos85_49 in85 sp49 3183.098862
Rwpos85_50 in85 sp50 3183.098862
Rwpos85_51 in85 sp51 3183.098862
Rwpos85_52 in85 sp52 3183.098862
Rwpos85_53 in85 sp53 3183.098862
Rwpos85_54 in85 sp54 3183.098862
Rwpos85_55 in85 sp55 11140.846016
Rwpos85_56 in85 sp56 3183.098862
Rwpos85_57 in85 sp57 3183.098862
Rwpos85_58 in85 sp58 3183.098862
Rwpos85_59 in85 sp59 11140.846016
Rwpos85_60 in85 sp60 11140.846016
Rwpos85_61 in85 sp61 11140.846016
Rwpos85_62 in85 sp62 11140.846016
Rwpos85_63 in85 sp63 3183.098862
Rwpos85_64 in85 sp64 11140.846016
Rwpos85_65 in85 sp65 3183.098862
Rwpos85_66 in85 sp66 3183.098862
Rwpos85_67 in85 sp67 3183.098862
Rwpos85_68 in85 sp68 3183.098862
Rwpos85_69 in85 sp69 3183.098862
Rwpos85_70 in85 sp70 3183.098862
Rwpos85_71 in85 sp71 3183.098862
Rwpos85_72 in85 sp72 11140.846016
Rwpos85_73 in85 sp73 11140.846016
Rwpos85_74 in85 sp74 11140.846016
Rwpos85_75 in85 sp75 11140.846016
Rwpos85_76 in85 sp76 11140.846016
Rwpos85_77 in85 sp77 11140.846016
Rwpos85_78 in85 sp78 3183.098862
Rwpos85_79 in85 sp79 3183.098862
Rwpos85_80 in85 sp80 11140.846016
Rwpos85_81 in85 sp81 3183.098862
Rwpos85_82 in85 sp82 3183.098862
Rwpos85_83 in85 sp83 3183.098862
Rwpos85_84 in85 sp84 11140.846016
Rwpos85_85 in85 sp85 3183.098862
Rwpos85_86 in85 sp86 11140.846016
Rwpos85_87 in85 sp87 11140.846016
Rwpos85_88 in85 sp88 3183.098862
Rwpos85_89 in85 sp89 11140.846016
Rwpos85_90 in85 sp90 3183.098862
Rwpos85_91 in85 sp91 11140.846016
Rwpos85_92 in85 sp92 3183.098862
Rwpos85_93 in85 sp93 3183.098862
Rwpos85_94 in85 sp94 11140.846016
Rwpos85_95 in85 sp95 11140.846016
Rwpos85_96 in85 sp96 3183.098862
Rwpos85_97 in85 sp97 3183.098862
Rwpos85_98 in85 sp98 3183.098862
Rwpos85_99 in85 sp99 3183.098862
Rwpos85_100 in85 sp100 3183.098862
Rwpos86_1 in86 sp1 3183.098862
Rwpos86_2 in86 sp2 11140.846016
Rwpos86_3 in86 sp3 3183.098862
Rwpos86_4 in86 sp4 11140.846016
Rwpos86_5 in86 sp5 3183.098862
Rwpos86_6 in86 sp6 3183.098862
Rwpos86_7 in86 sp7 3183.098862
Rwpos86_8 in86 sp8 3183.098862
Rwpos86_9 in86 sp9 11140.846016
Rwpos86_10 in86 sp10 3183.098862
Rwpos86_11 in86 sp11 3183.098862
Rwpos86_12 in86 sp12 11140.846016
Rwpos86_13 in86 sp13 3183.098862
Rwpos86_14 in86 sp14 3183.098862
Rwpos86_15 in86 sp15 11140.846016
Rwpos86_16 in86 sp16 3183.098862
Rwpos86_17 in86 sp17 3183.098862
Rwpos86_18 in86 sp18 11140.846016
Rwpos86_19 in86 sp19 3183.098862
Rwpos86_20 in86 sp20 3183.098862
Rwpos86_21 in86 sp21 11140.846016
Rwpos86_22 in86 sp22 3183.098862
Rwpos86_23 in86 sp23 3183.098862
Rwpos86_24 in86 sp24 11140.846016
Rwpos86_25 in86 sp25 3183.098862
Rwpos86_26 in86 sp26 11140.846016
Rwpos86_27 in86 sp27 3183.098862
Rwpos86_28 in86 sp28 3183.098862
Rwpos86_29 in86 sp29 11140.846016
Rwpos86_30 in86 sp30 3183.098862
Rwpos86_31 in86 sp31 11140.846016
Rwpos86_32 in86 sp32 3183.098862
Rwpos86_33 in86 sp33 3183.098862
Rwpos86_34 in86 sp34 11140.846016
Rwpos86_35 in86 sp35 11140.846016
Rwpos86_36 in86 sp36 11140.846016
Rwpos86_37 in86 sp37 3183.098862
Rwpos86_38 in86 sp38 3183.098862
Rwpos86_39 in86 sp39 11140.846016
Rwpos86_40 in86 sp40 11140.846016
Rwpos86_41 in86 sp41 11140.846016
Rwpos86_42 in86 sp42 11140.846016
Rwpos86_43 in86 sp43 11140.846016
Rwpos86_44 in86 sp44 11140.846016
Rwpos86_45 in86 sp45 11140.846016
Rwpos86_46 in86 sp46 11140.846016
Rwpos86_47 in86 sp47 3183.098862
Rwpos86_48 in86 sp48 11140.846016
Rwpos86_49 in86 sp49 11140.846016
Rwpos86_50 in86 sp50 11140.846016
Rwpos86_51 in86 sp51 11140.846016
Rwpos86_52 in86 sp52 3183.098862
Rwpos86_53 in86 sp53 11140.846016
Rwpos86_54 in86 sp54 11140.846016
Rwpos86_55 in86 sp55 3183.098862
Rwpos86_56 in86 sp56 3183.098862
Rwpos86_57 in86 sp57 3183.098862
Rwpos86_58 in86 sp58 3183.098862
Rwpos86_59 in86 sp59 11140.846016
Rwpos86_60 in86 sp60 11140.846016
Rwpos86_61 in86 sp61 11140.846016
Rwpos86_62 in86 sp62 11140.846016
Rwpos86_63 in86 sp63 11140.846016
Rwpos86_64 in86 sp64 3183.098862
Rwpos86_65 in86 sp65 3183.098862
Rwpos86_66 in86 sp66 11140.846016
Rwpos86_67 in86 sp67 3183.098862
Rwpos86_68 in86 sp68 3183.098862
Rwpos86_69 in86 sp69 11140.846016
Rwpos86_70 in86 sp70 11140.846016
Rwpos86_71 in86 sp71 11140.846016
Rwpos86_72 in86 sp72 11140.846016
Rwpos86_73 in86 sp73 3183.098862
Rwpos86_74 in86 sp74 11140.846016
Rwpos86_75 in86 sp75 3183.098862
Rwpos86_76 in86 sp76 3183.098862
Rwpos86_77 in86 sp77 11140.846016
Rwpos86_78 in86 sp78 3183.098862
Rwpos86_79 in86 sp79 3183.098862
Rwpos86_80 in86 sp80 3183.098862
Rwpos86_81 in86 sp81 11140.846016
Rwpos86_82 in86 sp82 11140.846016
Rwpos86_83 in86 sp83 3183.098862
Rwpos86_84 in86 sp84 3183.098862
Rwpos86_85 in86 sp85 11140.846016
Rwpos86_86 in86 sp86 3183.098862
Rwpos86_87 in86 sp87 11140.846016
Rwpos86_88 in86 sp88 3183.098862
Rwpos86_89 in86 sp89 11140.846016
Rwpos86_90 in86 sp90 3183.098862
Rwpos86_91 in86 sp91 3183.098862
Rwpos86_92 in86 sp92 11140.846016
Rwpos86_93 in86 sp93 11140.846016
Rwpos86_94 in86 sp94 3183.098862
Rwpos86_95 in86 sp95 3183.098862
Rwpos86_96 in86 sp96 3183.098862
Rwpos86_97 in86 sp97 3183.098862
Rwpos86_98 in86 sp98 11140.846016
Rwpos86_99 in86 sp99 11140.846016
Rwpos86_100 in86 sp100 3183.098862
Rwpos87_1 in87 sp1 3183.098862
Rwpos87_2 in87 sp2 3183.098862
Rwpos87_3 in87 sp3 11140.846016
Rwpos87_4 in87 sp4 11140.846016
Rwpos87_5 in87 sp5 11140.846016
Rwpos87_6 in87 sp6 3183.098862
Rwpos87_7 in87 sp7 3183.098862
Rwpos87_8 in87 sp8 11140.846016
Rwpos87_9 in87 sp9 3183.098862
Rwpos87_10 in87 sp10 3183.098862
Rwpos87_11 in87 sp11 3183.098862
Rwpos87_12 in87 sp12 3183.098862
Rwpos87_13 in87 sp13 11140.846016
Rwpos87_14 in87 sp14 3183.098862
Rwpos87_15 in87 sp15 11140.846016
Rwpos87_16 in87 sp16 3183.098862
Rwpos87_17 in87 sp17 11140.846016
Rwpos87_18 in87 sp18 3183.098862
Rwpos87_19 in87 sp19 11140.846016
Rwpos87_20 in87 sp20 11140.846016
Rwpos87_21 in87 sp21 11140.846016
Rwpos87_22 in87 sp22 3183.098862
Rwpos87_23 in87 sp23 3183.098862
Rwpos87_24 in87 sp24 3183.098862
Rwpos87_25 in87 sp25 3183.098862
Rwpos87_26 in87 sp26 3183.098862
Rwpos87_27 in87 sp27 3183.098862
Rwpos87_28 in87 sp28 3183.098862
Rwpos87_29 in87 sp29 11140.846016
Rwpos87_30 in87 sp30 3183.098862
Rwpos87_31 in87 sp31 3183.098862
Rwpos87_32 in87 sp32 3183.098862
Rwpos87_33 in87 sp33 3183.098862
Rwpos87_34 in87 sp34 3183.098862
Rwpos87_35 in87 sp35 3183.098862
Rwpos87_36 in87 sp36 11140.846016
Rwpos87_37 in87 sp37 11140.846016
Rwpos87_38 in87 sp38 11140.846016
Rwpos87_39 in87 sp39 3183.098862
Rwpos87_40 in87 sp40 11140.846016
Rwpos87_41 in87 sp41 3183.098862
Rwpos87_42 in87 sp42 11140.846016
Rwpos87_43 in87 sp43 3183.098862
Rwpos87_44 in87 sp44 3183.098862
Rwpos87_45 in87 sp45 3183.098862
Rwpos87_46 in87 sp46 3183.098862
Rwpos87_47 in87 sp47 11140.846016
Rwpos87_48 in87 sp48 3183.098862
Rwpos87_49 in87 sp49 11140.846016
Rwpos87_50 in87 sp50 3183.098862
Rwpos87_51 in87 sp51 11140.846016
Rwpos87_52 in87 sp52 3183.098862
Rwpos87_53 in87 sp53 11140.846016
Rwpos87_54 in87 sp54 11140.846016
Rwpos87_55 in87 sp55 11140.846016
Rwpos87_56 in87 sp56 11140.846016
Rwpos87_57 in87 sp57 3183.098862
Rwpos87_58 in87 sp58 11140.846016
Rwpos87_59 in87 sp59 3183.098862
Rwpos87_60 in87 sp60 11140.846016
Rwpos87_61 in87 sp61 11140.846016
Rwpos87_62 in87 sp62 3183.098862
Rwpos87_63 in87 sp63 11140.846016
Rwpos87_64 in87 sp64 3183.098862
Rwpos87_65 in87 sp65 11140.846016
Rwpos87_66 in87 sp66 11140.846016
Rwpos87_67 in87 sp67 3183.098862
Rwpos87_68 in87 sp68 11140.846016
Rwpos87_69 in87 sp69 11140.846016
Rwpos87_70 in87 sp70 11140.846016
Rwpos87_71 in87 sp71 11140.846016
Rwpos87_72 in87 sp72 11140.846016
Rwpos87_73 in87 sp73 3183.098862
Rwpos87_74 in87 sp74 11140.846016
Rwpos87_75 in87 sp75 3183.098862
Rwpos87_76 in87 sp76 3183.098862
Rwpos87_77 in87 sp77 11140.846016
Rwpos87_78 in87 sp78 11140.846016
Rwpos87_79 in87 sp79 11140.846016
Rwpos87_80 in87 sp80 3183.098862
Rwpos87_81 in87 sp81 3183.098862
Rwpos87_82 in87 sp82 11140.846016
Rwpos87_83 in87 sp83 3183.098862
Rwpos87_84 in87 sp84 11140.846016
Rwpos87_85 in87 sp85 11140.846016
Rwpos87_86 in87 sp86 11140.846016
Rwpos87_87 in87 sp87 11140.846016
Rwpos87_88 in87 sp88 11140.846016
Rwpos87_89 in87 sp89 3183.098862
Rwpos87_90 in87 sp90 11140.846016
Rwpos87_91 in87 sp91 3183.098862
Rwpos87_92 in87 sp92 3183.098862
Rwpos87_93 in87 sp93 3183.098862
Rwpos87_94 in87 sp94 11140.846016
Rwpos87_95 in87 sp95 3183.098862
Rwpos87_96 in87 sp96 3183.098862
Rwpos87_97 in87 sp97 3183.098862
Rwpos87_98 in87 sp98 11140.846016
Rwpos87_99 in87 sp99 3183.098862
Rwpos87_100 in87 sp100 11140.846016
Rwpos88_1 in88 sp1 3183.098862
Rwpos88_2 in88 sp2 11140.846016
Rwpos88_3 in88 sp3 11140.846016
Rwpos88_4 in88 sp4 11140.846016
Rwpos88_5 in88 sp5 3183.098862
Rwpos88_6 in88 sp6 3183.098862
Rwpos88_7 in88 sp7 3183.098862
Rwpos88_8 in88 sp8 11140.846016
Rwpos88_9 in88 sp9 11140.846016
Rwpos88_10 in88 sp10 11140.846016
Rwpos88_11 in88 sp11 3183.098862
Rwpos88_12 in88 sp12 3183.098862
Rwpos88_13 in88 sp13 3183.098862
Rwpos88_14 in88 sp14 3183.098862
Rwpos88_15 in88 sp15 3183.098862
Rwpos88_16 in88 sp16 11140.846016
Rwpos88_17 in88 sp17 11140.846016
Rwpos88_18 in88 sp18 11140.846016
Rwpos88_19 in88 sp19 3183.098862
Rwpos88_20 in88 sp20 11140.846016
Rwpos88_21 in88 sp21 3183.098862
Rwpos88_22 in88 sp22 3183.098862
Rwpos88_23 in88 sp23 3183.098862
Rwpos88_24 in88 sp24 11140.846016
Rwpos88_25 in88 sp25 11140.846016
Rwpos88_26 in88 sp26 3183.098862
Rwpos88_27 in88 sp27 11140.846016
Rwpos88_28 in88 sp28 3183.098862
Rwpos88_29 in88 sp29 3183.098862
Rwpos88_30 in88 sp30 11140.846016
Rwpos88_31 in88 sp31 11140.846016
Rwpos88_32 in88 sp32 11140.846016
Rwpos88_33 in88 sp33 3183.098862
Rwpos88_34 in88 sp34 3183.098862
Rwpos88_35 in88 sp35 11140.846016
Rwpos88_36 in88 sp36 11140.846016
Rwpos88_37 in88 sp37 3183.098862
Rwpos88_38 in88 sp38 3183.098862
Rwpos88_39 in88 sp39 3183.098862
Rwpos88_40 in88 sp40 3183.098862
Rwpos88_41 in88 sp41 11140.846016
Rwpos88_42 in88 sp42 3183.098862
Rwpos88_43 in88 sp43 11140.846016
Rwpos88_44 in88 sp44 3183.098862
Rwpos88_45 in88 sp45 11140.846016
Rwpos88_46 in88 sp46 3183.098862
Rwpos88_47 in88 sp47 3183.098862
Rwpos88_48 in88 sp48 11140.846016
Rwpos88_49 in88 sp49 3183.098862
Rwpos88_50 in88 sp50 3183.098862
Rwpos88_51 in88 sp51 3183.098862
Rwpos88_52 in88 sp52 11140.846016
Rwpos88_53 in88 sp53 3183.098862
Rwpos88_54 in88 sp54 3183.098862
Rwpos88_55 in88 sp55 3183.098862
Rwpos88_56 in88 sp56 11140.846016
Rwpos88_57 in88 sp57 11140.846016
Rwpos88_58 in88 sp58 3183.098862
Rwpos88_59 in88 sp59 11140.846016
Rwpos88_60 in88 sp60 11140.846016
Rwpos88_61 in88 sp61 3183.098862
Rwpos88_62 in88 sp62 11140.846016
Rwpos88_63 in88 sp63 3183.098862
Rwpos88_64 in88 sp64 3183.098862
Rwpos88_65 in88 sp65 11140.846016
Rwpos88_66 in88 sp66 3183.098862
Rwpos88_67 in88 sp67 3183.098862
Rwpos88_68 in88 sp68 11140.846016
Rwpos88_69 in88 sp69 11140.846016
Rwpos88_70 in88 sp70 3183.098862
Rwpos88_71 in88 sp71 3183.098862
Rwpos88_72 in88 sp72 3183.098862
Rwpos88_73 in88 sp73 11140.846016
Rwpos88_74 in88 sp74 11140.846016
Rwpos88_75 in88 sp75 3183.098862
Rwpos88_76 in88 sp76 3183.098862
Rwpos88_77 in88 sp77 11140.846016
Rwpos88_78 in88 sp78 3183.098862
Rwpos88_79 in88 sp79 11140.846016
Rwpos88_80 in88 sp80 11140.846016
Rwpos88_81 in88 sp81 11140.846016
Rwpos88_82 in88 sp82 3183.098862
Rwpos88_83 in88 sp83 11140.846016
Rwpos88_84 in88 sp84 11140.846016
Rwpos88_85 in88 sp85 11140.846016
Rwpos88_86 in88 sp86 3183.098862
Rwpos88_87 in88 sp87 3183.098862
Rwpos88_88 in88 sp88 3183.098862
Rwpos88_89 in88 sp89 3183.098862
Rwpos88_90 in88 sp90 11140.846016
Rwpos88_91 in88 sp91 11140.846016
Rwpos88_92 in88 sp92 11140.846016
Rwpos88_93 in88 sp93 3183.098862
Rwpos88_94 in88 sp94 11140.846016
Rwpos88_95 in88 sp95 11140.846016
Rwpos88_96 in88 sp96 11140.846016
Rwpos88_97 in88 sp97 3183.098862
Rwpos88_98 in88 sp98 11140.846016
Rwpos88_99 in88 sp99 3183.098862
Rwpos88_100 in88 sp100 3183.098862
Rwpos89_1 in89 sp1 3183.098862
Rwpos89_2 in89 sp2 3183.098862
Rwpos89_3 in89 sp3 3183.098862
Rwpos89_4 in89 sp4 3183.098862
Rwpos89_5 in89 sp5 11140.846016
Rwpos89_6 in89 sp6 11140.846016
Rwpos89_7 in89 sp7 11140.846016
Rwpos89_8 in89 sp8 3183.098862
Rwpos89_9 in89 sp9 3183.098862
Rwpos89_10 in89 sp10 11140.846016
Rwpos89_11 in89 sp11 11140.846016
Rwpos89_12 in89 sp12 3183.098862
Rwpos89_13 in89 sp13 3183.098862
Rwpos89_14 in89 sp14 3183.098862
Rwpos89_15 in89 sp15 3183.098862
Rwpos89_16 in89 sp16 11140.846016
Rwpos89_17 in89 sp17 11140.846016
Rwpos89_18 in89 sp18 3183.098862
Rwpos89_19 in89 sp19 3183.098862
Rwpos89_20 in89 sp20 3183.098862
Rwpos89_21 in89 sp21 11140.846016
Rwpos89_22 in89 sp22 11140.846016
Rwpos89_23 in89 sp23 3183.098862
Rwpos89_24 in89 sp24 3183.098862
Rwpos89_25 in89 sp25 11140.846016
Rwpos89_26 in89 sp26 11140.846016
Rwpos89_27 in89 sp27 11140.846016
Rwpos89_28 in89 sp28 11140.846016
Rwpos89_29 in89 sp29 11140.846016
Rwpos89_30 in89 sp30 3183.098862
Rwpos89_31 in89 sp31 3183.098862
Rwpos89_32 in89 sp32 3183.098862
Rwpos89_33 in89 sp33 11140.846016
Rwpos89_34 in89 sp34 3183.098862
Rwpos89_35 in89 sp35 11140.846016
Rwpos89_36 in89 sp36 3183.098862
Rwpos89_37 in89 sp37 11140.846016
Rwpos89_38 in89 sp38 11140.846016
Rwpos89_39 in89 sp39 11140.846016
Rwpos89_40 in89 sp40 3183.098862
Rwpos89_41 in89 sp41 3183.098862
Rwpos89_42 in89 sp42 3183.098862
Rwpos89_43 in89 sp43 11140.846016
Rwpos89_44 in89 sp44 3183.098862
Rwpos89_45 in89 sp45 3183.098862
Rwpos89_46 in89 sp46 11140.846016
Rwpos89_47 in89 sp47 3183.098862
Rwpos89_48 in89 sp48 11140.846016
Rwpos89_49 in89 sp49 3183.098862
Rwpos89_50 in89 sp50 3183.098862
Rwpos89_51 in89 sp51 3183.098862
Rwpos89_52 in89 sp52 3183.098862
Rwpos89_53 in89 sp53 11140.846016
Rwpos89_54 in89 sp54 11140.846016
Rwpos89_55 in89 sp55 11140.846016
Rwpos89_56 in89 sp56 3183.098862
Rwpos89_57 in89 sp57 3183.098862
Rwpos89_58 in89 sp58 3183.098862
Rwpos89_59 in89 sp59 11140.846016
Rwpos89_60 in89 sp60 11140.846016
Rwpos89_61 in89 sp61 11140.846016
Rwpos89_62 in89 sp62 3183.098862
Rwpos89_63 in89 sp63 3183.098862
Rwpos89_64 in89 sp64 11140.846016
Rwpos89_65 in89 sp65 11140.846016
Rwpos89_66 in89 sp66 3183.098862
Rwpos89_67 in89 sp67 11140.846016
Rwpos89_68 in89 sp68 3183.098862
Rwpos89_69 in89 sp69 3183.098862
Rwpos89_70 in89 sp70 3183.098862
Rwpos89_71 in89 sp71 3183.098862
Rwpos89_72 in89 sp72 3183.098862
Rwpos89_73 in89 sp73 11140.846016
Rwpos89_74 in89 sp74 3183.098862
Rwpos89_75 in89 sp75 11140.846016
Rwpos89_76 in89 sp76 11140.846016
Rwpos89_77 in89 sp77 11140.846016
Rwpos89_78 in89 sp78 3183.098862
Rwpos89_79 in89 sp79 3183.098862
Rwpos89_80 in89 sp80 11140.846016
Rwpos89_81 in89 sp81 11140.846016
Rwpos89_82 in89 sp82 3183.098862
Rwpos89_83 in89 sp83 3183.098862
Rwpos89_84 in89 sp84 3183.098862
Rwpos89_85 in89 sp85 3183.098862
Rwpos89_86 in89 sp86 3183.098862
Rwpos89_87 in89 sp87 3183.098862
Rwpos89_88 in89 sp88 3183.098862
Rwpos89_89 in89 sp89 11140.846016
Rwpos89_90 in89 sp90 3183.098862
Rwpos89_91 in89 sp91 11140.846016
Rwpos89_92 in89 sp92 11140.846016
Rwpos89_93 in89 sp93 3183.098862
Rwpos89_94 in89 sp94 11140.846016
Rwpos89_95 in89 sp95 3183.098862
Rwpos89_96 in89 sp96 11140.846016
Rwpos89_97 in89 sp97 3183.098862
Rwpos89_98 in89 sp98 3183.098862
Rwpos89_99 in89 sp99 3183.098862
Rwpos89_100 in89 sp100 11140.846016
Rwpos90_1 in90 sp1 3183.098862
Rwpos90_2 in90 sp2 3183.098862
Rwpos90_3 in90 sp3 3183.098862
Rwpos90_4 in90 sp4 11140.846016
Rwpos90_5 in90 sp5 11140.846016
Rwpos90_6 in90 sp6 3183.098862
Rwpos90_7 in90 sp7 11140.846016
Rwpos90_8 in90 sp8 11140.846016
Rwpos90_9 in90 sp9 11140.846016
Rwpos90_10 in90 sp10 3183.098862
Rwpos90_11 in90 sp11 11140.846016
Rwpos90_12 in90 sp12 11140.846016
Rwpos90_13 in90 sp13 11140.846016
Rwpos90_14 in90 sp14 3183.098862
Rwpos90_15 in90 sp15 3183.098862
Rwpos90_16 in90 sp16 11140.846016
Rwpos90_17 in90 sp17 11140.846016
Rwpos90_18 in90 sp18 3183.098862
Rwpos90_19 in90 sp19 3183.098862
Rwpos90_20 in90 sp20 3183.098862
Rwpos90_21 in90 sp21 11140.846016
Rwpos90_22 in90 sp22 3183.098862
Rwpos90_23 in90 sp23 11140.846016
Rwpos90_24 in90 sp24 3183.098862
Rwpos90_25 in90 sp25 3183.098862
Rwpos90_26 in90 sp26 3183.098862
Rwpos90_27 in90 sp27 11140.846016
Rwpos90_28 in90 sp28 11140.846016
Rwpos90_29 in90 sp29 11140.846016
Rwpos90_30 in90 sp30 11140.846016
Rwpos90_31 in90 sp31 11140.846016
Rwpos90_32 in90 sp32 11140.846016
Rwpos90_33 in90 sp33 11140.846016
Rwpos90_34 in90 sp34 3183.098862
Rwpos90_35 in90 sp35 3183.098862
Rwpos90_36 in90 sp36 3183.098862
Rwpos90_37 in90 sp37 11140.846016
Rwpos90_38 in90 sp38 11140.846016
Rwpos90_39 in90 sp39 11140.846016
Rwpos90_40 in90 sp40 11140.846016
Rwpos90_41 in90 sp41 11140.846016
Rwpos90_42 in90 sp42 3183.098862
Rwpos90_43 in90 sp43 11140.846016
Rwpos90_44 in90 sp44 11140.846016
Rwpos90_45 in90 sp45 11140.846016
Rwpos90_46 in90 sp46 11140.846016
Rwpos90_47 in90 sp47 11140.846016
Rwpos90_48 in90 sp48 3183.098862
Rwpos90_49 in90 sp49 3183.098862
Rwpos90_50 in90 sp50 3183.098862
Rwpos90_51 in90 sp51 11140.846016
Rwpos90_52 in90 sp52 3183.098862
Rwpos90_53 in90 sp53 11140.846016
Rwpos90_54 in90 sp54 11140.846016
Rwpos90_55 in90 sp55 3183.098862
Rwpos90_56 in90 sp56 11140.846016
Rwpos90_57 in90 sp57 11140.846016
Rwpos90_58 in90 sp58 11140.846016
Rwpos90_59 in90 sp59 11140.846016
Rwpos90_60 in90 sp60 11140.846016
Rwpos90_61 in90 sp61 11140.846016
Rwpos90_62 in90 sp62 3183.098862
Rwpos90_63 in90 sp63 11140.846016
Rwpos90_64 in90 sp64 3183.098862
Rwpos90_65 in90 sp65 11140.846016
Rwpos90_66 in90 sp66 11140.846016
Rwpos90_67 in90 sp67 3183.098862
Rwpos90_68 in90 sp68 3183.098862
Rwpos90_69 in90 sp69 11140.846016
Rwpos90_70 in90 sp70 11140.846016
Rwpos90_71 in90 sp71 11140.846016
Rwpos90_72 in90 sp72 11140.846016
Rwpos90_73 in90 sp73 11140.846016
Rwpos90_74 in90 sp74 11140.846016
Rwpos90_75 in90 sp75 3183.098862
Rwpos90_76 in90 sp76 11140.846016
Rwpos90_77 in90 sp77 3183.098862
Rwpos90_78 in90 sp78 11140.846016
Rwpos90_79 in90 sp79 11140.846016
Rwpos90_80 in90 sp80 11140.846016
Rwpos90_81 in90 sp81 3183.098862
Rwpos90_82 in90 sp82 11140.846016
Rwpos90_83 in90 sp83 11140.846016
Rwpos90_84 in90 sp84 11140.846016
Rwpos90_85 in90 sp85 3183.098862
Rwpos90_86 in90 sp86 11140.846016
Rwpos90_87 in90 sp87 3183.098862
Rwpos90_88 in90 sp88 11140.846016
Rwpos90_89 in90 sp89 11140.846016
Rwpos90_90 in90 sp90 11140.846016
Rwpos90_91 in90 sp91 11140.846016
Rwpos90_92 in90 sp92 3183.098862
Rwpos90_93 in90 sp93 11140.846016
Rwpos90_94 in90 sp94 3183.098862
Rwpos90_95 in90 sp95 3183.098862
Rwpos90_96 in90 sp96 11140.846016
Rwpos90_97 in90 sp97 3183.098862
Rwpos90_98 in90 sp98 3183.098862
Rwpos90_99 in90 sp99 11140.846016
Rwpos90_100 in90 sp100 3183.098862
Rwpos91_1 in91 sp1 11140.846016
Rwpos91_2 in91 sp2 11140.846016
Rwpos91_3 in91 sp3 11140.846016
Rwpos91_4 in91 sp4 3183.098862
Rwpos91_5 in91 sp5 11140.846016
Rwpos91_6 in91 sp6 3183.098862
Rwpos91_7 in91 sp7 11140.846016
Rwpos91_8 in91 sp8 3183.098862
Rwpos91_9 in91 sp9 11140.846016
Rwpos91_10 in91 sp10 11140.846016
Rwpos91_11 in91 sp11 11140.846016
Rwpos91_12 in91 sp12 11140.846016
Rwpos91_13 in91 sp13 11140.846016
Rwpos91_14 in91 sp14 11140.846016
Rwpos91_15 in91 sp15 3183.098862
Rwpos91_16 in91 sp16 3183.098862
Rwpos91_17 in91 sp17 11140.846016
Rwpos91_18 in91 sp18 11140.846016
Rwpos91_19 in91 sp19 11140.846016
Rwpos91_20 in91 sp20 3183.098862
Rwpos91_21 in91 sp21 3183.098862
Rwpos91_22 in91 sp22 3183.098862
Rwpos91_23 in91 sp23 3183.098862
Rwpos91_24 in91 sp24 11140.846016
Rwpos91_25 in91 sp25 11140.846016
Rwpos91_26 in91 sp26 3183.098862
Rwpos91_27 in91 sp27 11140.846016
Rwpos91_28 in91 sp28 3183.098862
Rwpos91_29 in91 sp29 3183.098862
Rwpos91_30 in91 sp30 11140.846016
Rwpos91_31 in91 sp31 11140.846016
Rwpos91_32 in91 sp32 3183.098862
Rwpos91_33 in91 sp33 3183.098862
Rwpos91_34 in91 sp34 3183.098862
Rwpos91_35 in91 sp35 11140.846016
Rwpos91_36 in91 sp36 3183.098862
Rwpos91_37 in91 sp37 3183.098862
Rwpos91_38 in91 sp38 11140.846016
Rwpos91_39 in91 sp39 11140.846016
Rwpos91_40 in91 sp40 11140.846016
Rwpos91_41 in91 sp41 11140.846016
Rwpos91_42 in91 sp42 3183.098862
Rwpos91_43 in91 sp43 3183.098862
Rwpos91_44 in91 sp44 3183.098862
Rwpos91_45 in91 sp45 11140.846016
Rwpos91_46 in91 sp46 3183.098862
Rwpos91_47 in91 sp47 3183.098862
Rwpos91_48 in91 sp48 11140.846016
Rwpos91_49 in91 sp49 3183.098862
Rwpos91_50 in91 sp50 3183.098862
Rwpos91_51 in91 sp51 11140.846016
Rwpos91_52 in91 sp52 11140.846016
Rwpos91_53 in91 sp53 11140.846016
Rwpos91_54 in91 sp54 3183.098862
Rwpos91_55 in91 sp55 3183.098862
Rwpos91_56 in91 sp56 3183.098862
Rwpos91_57 in91 sp57 3183.098862
Rwpos91_58 in91 sp58 3183.098862
Rwpos91_59 in91 sp59 3183.098862
Rwpos91_60 in91 sp60 3183.098862
Rwpos91_61 in91 sp61 11140.846016
Rwpos91_62 in91 sp62 3183.098862
Rwpos91_63 in91 sp63 11140.846016
Rwpos91_64 in91 sp64 3183.098862
Rwpos91_65 in91 sp65 11140.846016
Rwpos91_66 in91 sp66 3183.098862
Rwpos91_67 in91 sp67 11140.846016
Rwpos91_68 in91 sp68 11140.846016
Rwpos91_69 in91 sp69 11140.846016
Rwpos91_70 in91 sp70 3183.098862
Rwpos91_71 in91 sp71 11140.846016
Rwpos91_72 in91 sp72 11140.846016
Rwpos91_73 in91 sp73 11140.846016
Rwpos91_74 in91 sp74 11140.846016
Rwpos91_75 in91 sp75 3183.098862
Rwpos91_76 in91 sp76 3183.098862
Rwpos91_77 in91 sp77 3183.098862
Rwpos91_78 in91 sp78 3183.098862
Rwpos91_79 in91 sp79 11140.846016
Rwpos91_80 in91 sp80 3183.098862
Rwpos91_81 in91 sp81 11140.846016
Rwpos91_82 in91 sp82 3183.098862
Rwpos91_83 in91 sp83 11140.846016
Rwpos91_84 in91 sp84 3183.098862
Rwpos91_85 in91 sp85 11140.846016
Rwpos91_86 in91 sp86 3183.098862
Rwpos91_87 in91 sp87 3183.098862
Rwpos91_88 in91 sp88 11140.846016
Rwpos91_89 in91 sp89 3183.098862
Rwpos91_90 in91 sp90 11140.846016
Rwpos91_91 in91 sp91 3183.098862
Rwpos91_92 in91 sp92 3183.098862
Rwpos91_93 in91 sp93 11140.846016
Rwpos91_94 in91 sp94 3183.098862
Rwpos91_95 in91 sp95 11140.846016
Rwpos91_96 in91 sp96 3183.098862
Rwpos91_97 in91 sp97 11140.846016
Rwpos91_98 in91 sp98 3183.098862
Rwpos91_99 in91 sp99 11140.846016
Rwpos91_100 in91 sp100 11140.846016
Rwpos92_1 in92 sp1 11140.846016
Rwpos92_2 in92 sp2 11140.846016
Rwpos92_3 in92 sp3 3183.098862
Rwpos92_4 in92 sp4 11140.846016
Rwpos92_5 in92 sp5 3183.098862
Rwpos92_6 in92 sp6 3183.098862
Rwpos92_7 in92 sp7 3183.098862
Rwpos92_8 in92 sp8 3183.098862
Rwpos92_9 in92 sp9 11140.846016
Rwpos92_10 in92 sp10 11140.846016
Rwpos92_11 in92 sp11 3183.098862
Rwpos92_12 in92 sp12 3183.098862
Rwpos92_13 in92 sp13 11140.846016
Rwpos92_14 in92 sp14 3183.098862
Rwpos92_15 in92 sp15 3183.098862
Rwpos92_16 in92 sp16 11140.846016
Rwpos92_17 in92 sp17 3183.098862
Rwpos92_18 in92 sp18 11140.846016
Rwpos92_19 in92 sp19 3183.098862
Rwpos92_20 in92 sp20 11140.846016
Rwpos92_21 in92 sp21 3183.098862
Rwpos92_22 in92 sp22 3183.098862
Rwpos92_23 in92 sp23 3183.098862
Rwpos92_24 in92 sp24 11140.846016
Rwpos92_25 in92 sp25 3183.098862
Rwpos92_26 in92 sp26 3183.098862
Rwpos92_27 in92 sp27 3183.098862
Rwpos92_28 in92 sp28 3183.098862
Rwpos92_29 in92 sp29 11140.846016
Rwpos92_30 in92 sp30 3183.098862
Rwpos92_31 in92 sp31 11140.846016
Rwpos92_32 in92 sp32 11140.846016
Rwpos92_33 in92 sp33 11140.846016
Rwpos92_34 in92 sp34 11140.846016
Rwpos92_35 in92 sp35 3183.098862
Rwpos92_36 in92 sp36 11140.846016
Rwpos92_37 in92 sp37 3183.098862
Rwpos92_38 in92 sp38 3183.098862
Rwpos92_39 in92 sp39 3183.098862
Rwpos92_40 in92 sp40 11140.846016
Rwpos92_41 in92 sp41 3183.098862
Rwpos92_42 in92 sp42 11140.846016
Rwpos92_43 in92 sp43 11140.846016
Rwpos92_44 in92 sp44 3183.098862
Rwpos92_45 in92 sp45 11140.846016
Rwpos92_46 in92 sp46 11140.846016
Rwpos92_47 in92 sp47 3183.098862
Rwpos92_48 in92 sp48 11140.846016
Rwpos92_49 in92 sp49 11140.846016
Rwpos92_50 in92 sp50 3183.098862
Rwpos92_51 in92 sp51 11140.846016
Rwpos92_52 in92 sp52 11140.846016
Rwpos92_53 in92 sp53 11140.846016
Rwpos92_54 in92 sp54 3183.098862
Rwpos92_55 in92 sp55 3183.098862
Rwpos92_56 in92 sp56 11140.846016
Rwpos92_57 in92 sp57 3183.098862
Rwpos92_58 in92 sp58 11140.846016
Rwpos92_59 in92 sp59 11140.846016
Rwpos92_60 in92 sp60 3183.098862
Rwpos92_61 in92 sp61 11140.846016
Rwpos92_62 in92 sp62 11140.846016
Rwpos92_63 in92 sp63 3183.098862
Rwpos92_64 in92 sp64 11140.846016
Rwpos92_65 in92 sp65 11140.846016
Rwpos92_66 in92 sp66 11140.846016
Rwpos92_67 in92 sp67 11140.846016
Rwpos92_68 in92 sp68 11140.846016
Rwpos92_69 in92 sp69 3183.098862
Rwpos92_70 in92 sp70 3183.098862
Rwpos92_71 in92 sp71 3183.098862
Rwpos92_72 in92 sp72 11140.846016
Rwpos92_73 in92 sp73 11140.846016
Rwpos92_74 in92 sp74 11140.846016
Rwpos92_75 in92 sp75 3183.098862
Rwpos92_76 in92 sp76 3183.098862
Rwpos92_77 in92 sp77 11140.846016
Rwpos92_78 in92 sp78 11140.846016
Rwpos92_79 in92 sp79 3183.098862
Rwpos92_80 in92 sp80 3183.098862
Rwpos92_81 in92 sp81 3183.098862
Rwpos92_82 in92 sp82 3183.098862
Rwpos92_83 in92 sp83 11140.846016
Rwpos92_84 in92 sp84 3183.098862
Rwpos92_85 in92 sp85 3183.098862
Rwpos92_86 in92 sp86 3183.098862
Rwpos92_87 in92 sp87 3183.098862
Rwpos92_88 in92 sp88 11140.846016
Rwpos92_89 in92 sp89 11140.846016
Rwpos92_90 in92 sp90 11140.846016
Rwpos92_91 in92 sp91 11140.846016
Rwpos92_92 in92 sp92 3183.098862
Rwpos92_93 in92 sp93 3183.098862
Rwpos92_94 in92 sp94 11140.846016
Rwpos92_95 in92 sp95 3183.098862
Rwpos92_96 in92 sp96 3183.098862
Rwpos92_97 in92 sp97 11140.846016
Rwpos92_98 in92 sp98 3183.098862
Rwpos92_99 in92 sp99 11140.846016
Rwpos92_100 in92 sp100 11140.846016
Rwpos93_1 in93 sp1 3183.098862
Rwpos93_2 in93 sp2 3183.098862
Rwpos93_3 in93 sp3 3183.098862
Rwpos93_4 in93 sp4 3183.098862
Rwpos93_5 in93 sp5 3183.098862
Rwpos93_6 in93 sp6 11140.846016
Rwpos93_7 in93 sp7 3183.098862
Rwpos93_8 in93 sp8 3183.098862
Rwpos93_9 in93 sp9 11140.846016
Rwpos93_10 in93 sp10 11140.846016
Rwpos93_11 in93 sp11 11140.846016
Rwpos93_12 in93 sp12 3183.098862
Rwpos93_13 in93 sp13 3183.098862
Rwpos93_14 in93 sp14 3183.098862
Rwpos93_15 in93 sp15 3183.098862
Rwpos93_16 in93 sp16 11140.846016
Rwpos93_17 in93 sp17 3183.098862
Rwpos93_18 in93 sp18 3183.098862
Rwpos93_19 in93 sp19 3183.098862
Rwpos93_20 in93 sp20 3183.098862
Rwpos93_21 in93 sp21 3183.098862
Rwpos93_22 in93 sp22 3183.098862
Rwpos93_23 in93 sp23 3183.098862
Rwpos93_24 in93 sp24 3183.098862
Rwpos93_25 in93 sp25 3183.098862
Rwpos93_26 in93 sp26 11140.846016
Rwpos93_27 in93 sp27 11140.846016
Rwpos93_28 in93 sp28 3183.098862
Rwpos93_29 in93 sp29 3183.098862
Rwpos93_30 in93 sp30 11140.846016
Rwpos93_31 in93 sp31 3183.098862
Rwpos93_32 in93 sp32 11140.846016
Rwpos93_33 in93 sp33 11140.846016
Rwpos93_34 in93 sp34 3183.098862
Rwpos93_35 in93 sp35 3183.098862
Rwpos93_36 in93 sp36 3183.098862
Rwpos93_37 in93 sp37 3183.098862
Rwpos93_38 in93 sp38 11140.846016
Rwpos93_39 in93 sp39 11140.846016
Rwpos93_40 in93 sp40 3183.098862
Rwpos93_41 in93 sp41 11140.846016
Rwpos93_42 in93 sp42 11140.846016
Rwpos93_43 in93 sp43 3183.098862
Rwpos93_44 in93 sp44 11140.846016
Rwpos93_45 in93 sp45 3183.098862
Rwpos93_46 in93 sp46 3183.098862
Rwpos93_47 in93 sp47 3183.098862
Rwpos93_48 in93 sp48 11140.846016
Rwpos93_49 in93 sp49 3183.098862
Rwpos93_50 in93 sp50 3183.098862
Rwpos93_51 in93 sp51 3183.098862
Rwpos93_52 in93 sp52 3183.098862
Rwpos93_53 in93 sp53 3183.098862
Rwpos93_54 in93 sp54 11140.846016
Rwpos93_55 in93 sp55 11140.846016
Rwpos93_56 in93 sp56 3183.098862
Rwpos93_57 in93 sp57 3183.098862
Rwpos93_58 in93 sp58 3183.098862
Rwpos93_59 in93 sp59 11140.846016
Rwpos93_60 in93 sp60 3183.098862
Rwpos93_61 in93 sp61 11140.846016
Rwpos93_62 in93 sp62 11140.846016
Rwpos93_63 in93 sp63 3183.098862
Rwpos93_64 in93 sp64 11140.846016
Rwpos93_65 in93 sp65 3183.098862
Rwpos93_66 in93 sp66 3183.098862
Rwpos93_67 in93 sp67 3183.098862
Rwpos93_68 in93 sp68 3183.098862
Rwpos93_69 in93 sp69 3183.098862
Rwpos93_70 in93 sp70 3183.098862
Rwpos93_71 in93 sp71 11140.846016
Rwpos93_72 in93 sp72 3183.098862
Rwpos93_73 in93 sp73 3183.098862
Rwpos93_74 in93 sp74 3183.098862
Rwpos93_75 in93 sp75 11140.846016
Rwpos93_76 in93 sp76 3183.098862
Rwpos93_77 in93 sp77 3183.098862
Rwpos93_78 in93 sp78 3183.098862
Rwpos93_79 in93 sp79 3183.098862
Rwpos93_80 in93 sp80 11140.846016
Rwpos93_81 in93 sp81 3183.098862
Rwpos93_82 in93 sp82 3183.098862
Rwpos93_83 in93 sp83 3183.098862
Rwpos93_84 in93 sp84 3183.098862
Rwpos93_85 in93 sp85 3183.098862
Rwpos93_86 in93 sp86 11140.846016
Rwpos93_87 in93 sp87 3183.098862
Rwpos93_88 in93 sp88 3183.098862
Rwpos93_89 in93 sp89 11140.846016
Rwpos93_90 in93 sp90 11140.846016
Rwpos93_91 in93 sp91 11140.846016
Rwpos93_92 in93 sp92 11140.846016
Rwpos93_93 in93 sp93 11140.846016
Rwpos93_94 in93 sp94 11140.846016
Rwpos93_95 in93 sp95 3183.098862
Rwpos93_96 in93 sp96 11140.846016
Rwpos93_97 in93 sp97 11140.846016
Rwpos93_98 in93 sp98 3183.098862
Rwpos93_99 in93 sp99 3183.098862
Rwpos93_100 in93 sp100 3183.098862
Rwpos94_1 in94 sp1 3183.098862
Rwpos94_2 in94 sp2 11140.846016
Rwpos94_3 in94 sp3 3183.098862
Rwpos94_4 in94 sp4 3183.098862
Rwpos94_5 in94 sp5 3183.098862
Rwpos94_6 in94 sp6 3183.098862
Rwpos94_7 in94 sp7 3183.098862
Rwpos94_8 in94 sp8 11140.846016
Rwpos94_9 in94 sp9 11140.846016
Rwpos94_10 in94 sp10 11140.846016
Rwpos94_11 in94 sp11 3183.098862
Rwpos94_12 in94 sp12 3183.098862
Rwpos94_13 in94 sp13 3183.098862
Rwpos94_14 in94 sp14 11140.846016
Rwpos94_15 in94 sp15 11140.846016
Rwpos94_16 in94 sp16 3183.098862
Rwpos94_17 in94 sp17 3183.098862
Rwpos94_18 in94 sp18 3183.098862
Rwpos94_19 in94 sp19 3183.098862
Rwpos94_20 in94 sp20 3183.098862
Rwpos94_21 in94 sp21 11140.846016
Rwpos94_22 in94 sp22 3183.098862
Rwpos94_23 in94 sp23 11140.846016
Rwpos94_24 in94 sp24 3183.098862
Rwpos94_25 in94 sp25 11140.846016
Rwpos94_26 in94 sp26 11140.846016
Rwpos94_27 in94 sp27 3183.098862
Rwpos94_28 in94 sp28 11140.846016
Rwpos94_29 in94 sp29 11140.846016
Rwpos94_30 in94 sp30 3183.098862
Rwpos94_31 in94 sp31 3183.098862
Rwpos94_32 in94 sp32 3183.098862
Rwpos94_33 in94 sp33 11140.846016
Rwpos94_34 in94 sp34 3183.098862
Rwpos94_35 in94 sp35 3183.098862
Rwpos94_36 in94 sp36 3183.098862
Rwpos94_37 in94 sp37 3183.098862
Rwpos94_38 in94 sp38 3183.098862
Rwpos94_39 in94 sp39 11140.846016
Rwpos94_40 in94 sp40 11140.846016
Rwpos94_41 in94 sp41 3183.098862
Rwpos94_42 in94 sp42 11140.846016
Rwpos94_43 in94 sp43 3183.098862
Rwpos94_44 in94 sp44 11140.846016
Rwpos94_45 in94 sp45 3183.098862
Rwpos94_46 in94 sp46 3183.098862
Rwpos94_47 in94 sp47 3183.098862
Rwpos94_48 in94 sp48 11140.846016
Rwpos94_49 in94 sp49 11140.846016
Rwpos94_50 in94 sp50 3183.098862
Rwpos94_51 in94 sp51 11140.846016
Rwpos94_52 in94 sp52 11140.846016
Rwpos94_53 in94 sp53 3183.098862
Rwpos94_54 in94 sp54 3183.098862
Rwpos94_55 in94 sp55 11140.846016
Rwpos94_56 in94 sp56 11140.846016
Rwpos94_57 in94 sp57 3183.098862
Rwpos94_58 in94 sp58 11140.846016
Rwpos94_59 in94 sp59 3183.098862
Rwpos94_60 in94 sp60 3183.098862
Rwpos94_61 in94 sp61 3183.098862
Rwpos94_62 in94 sp62 3183.098862
Rwpos94_63 in94 sp63 11140.846016
Rwpos94_64 in94 sp64 11140.846016
Rwpos94_65 in94 sp65 11140.846016
Rwpos94_66 in94 sp66 11140.846016
Rwpos94_67 in94 sp67 11140.846016
Rwpos94_68 in94 sp68 3183.098862
Rwpos94_69 in94 sp69 11140.846016
Rwpos94_70 in94 sp70 11140.846016
Rwpos94_71 in94 sp71 3183.098862
Rwpos94_72 in94 sp72 11140.846016
Rwpos94_73 in94 sp73 3183.098862
Rwpos94_74 in94 sp74 11140.846016
Rwpos94_75 in94 sp75 11140.846016
Rwpos94_76 in94 sp76 3183.098862
Rwpos94_77 in94 sp77 3183.098862
Rwpos94_78 in94 sp78 3183.098862
Rwpos94_79 in94 sp79 11140.846016
Rwpos94_80 in94 sp80 11140.846016
Rwpos94_81 in94 sp81 11140.846016
Rwpos94_82 in94 sp82 11140.846016
Rwpos94_83 in94 sp83 3183.098862
Rwpos94_84 in94 sp84 11140.846016
Rwpos94_85 in94 sp85 3183.098862
Rwpos94_86 in94 sp86 3183.098862
Rwpos94_87 in94 sp87 11140.846016
Rwpos94_88 in94 sp88 11140.846016
Rwpos94_89 in94 sp89 11140.846016
Rwpos94_90 in94 sp90 3183.098862
Rwpos94_91 in94 sp91 11140.846016
Rwpos94_92 in94 sp92 3183.098862
Rwpos94_93 in94 sp93 3183.098862
Rwpos94_94 in94 sp94 3183.098862
Rwpos94_95 in94 sp95 3183.098862
Rwpos94_96 in94 sp96 3183.098862
Rwpos94_97 in94 sp97 3183.098862
Rwpos94_98 in94 sp98 3183.098862
Rwpos94_99 in94 sp99 3183.098862
Rwpos94_100 in94 sp100 3183.098862
Rwpos95_1 in95 sp1 11140.846016
Rwpos95_2 in95 sp2 3183.098862
Rwpos95_3 in95 sp3 11140.846016
Rwpos95_4 in95 sp4 11140.846016
Rwpos95_5 in95 sp5 11140.846016
Rwpos95_6 in95 sp6 3183.098862
Rwpos95_7 in95 sp7 11140.846016
Rwpos95_8 in95 sp8 3183.098862
Rwpos95_9 in95 sp9 3183.098862
Rwpos95_10 in95 sp10 3183.098862
Rwpos95_11 in95 sp11 3183.098862
Rwpos95_12 in95 sp12 11140.846016
Rwpos95_13 in95 sp13 11140.846016
Rwpos95_14 in95 sp14 3183.098862
Rwpos95_15 in95 sp15 3183.098862
Rwpos95_16 in95 sp16 11140.846016
Rwpos95_17 in95 sp17 3183.098862
Rwpos95_18 in95 sp18 3183.098862
Rwpos95_19 in95 sp19 11140.846016
Rwpos95_20 in95 sp20 3183.098862
Rwpos95_21 in95 sp21 3183.098862
Rwpos95_22 in95 sp22 3183.098862
Rwpos95_23 in95 sp23 3183.098862
Rwpos95_24 in95 sp24 3183.098862
Rwpos95_25 in95 sp25 11140.846016
Rwpos95_26 in95 sp26 3183.098862
Rwpos95_27 in95 sp27 3183.098862
Rwpos95_28 in95 sp28 3183.098862
Rwpos95_29 in95 sp29 3183.098862
Rwpos95_30 in95 sp30 11140.846016
Rwpos95_31 in95 sp31 3183.098862
Rwpos95_32 in95 sp32 3183.098862
Rwpos95_33 in95 sp33 11140.846016
Rwpos95_34 in95 sp34 3183.098862
Rwpos95_35 in95 sp35 3183.098862
Rwpos95_36 in95 sp36 11140.846016
Rwpos95_37 in95 sp37 3183.098862
Rwpos95_38 in95 sp38 3183.098862
Rwpos95_39 in95 sp39 3183.098862
Rwpos95_40 in95 sp40 3183.098862
Rwpos95_41 in95 sp41 11140.846016
Rwpos95_42 in95 sp42 3183.098862
Rwpos95_43 in95 sp43 3183.098862
Rwpos95_44 in95 sp44 11140.846016
Rwpos95_45 in95 sp45 3183.098862
Rwpos95_46 in95 sp46 11140.846016
Rwpos95_47 in95 sp47 3183.098862
Rwpos95_48 in95 sp48 11140.846016
Rwpos95_49 in95 sp49 11140.846016
Rwpos95_50 in95 sp50 11140.846016
Rwpos95_51 in95 sp51 11140.846016
Rwpos95_52 in95 sp52 11140.846016
Rwpos95_53 in95 sp53 3183.098862
Rwpos95_54 in95 sp54 3183.098862
Rwpos95_55 in95 sp55 3183.098862
Rwpos95_56 in95 sp56 11140.846016
Rwpos95_57 in95 sp57 11140.846016
Rwpos95_58 in95 sp58 11140.846016
Rwpos95_59 in95 sp59 3183.098862
Rwpos95_60 in95 sp60 11140.846016
Rwpos95_61 in95 sp61 3183.098862
Rwpos95_62 in95 sp62 11140.846016
Rwpos95_63 in95 sp63 3183.098862
Rwpos95_64 in95 sp64 11140.846016
Rwpos95_65 in95 sp65 11140.846016
Rwpos95_66 in95 sp66 3183.098862
Rwpos95_67 in95 sp67 11140.846016
Rwpos95_68 in95 sp68 3183.098862
Rwpos95_69 in95 sp69 3183.098862
Rwpos95_70 in95 sp70 3183.098862
Rwpos95_71 in95 sp71 3183.098862
Rwpos95_72 in95 sp72 3183.098862
Rwpos95_73 in95 sp73 3183.098862
Rwpos95_74 in95 sp74 3183.098862
Rwpos95_75 in95 sp75 3183.098862
Rwpos95_76 in95 sp76 3183.098862
Rwpos95_77 in95 sp77 11140.846016
Rwpos95_78 in95 sp78 11140.846016
Rwpos95_79 in95 sp79 11140.846016
Rwpos95_80 in95 sp80 3183.098862
Rwpos95_81 in95 sp81 3183.098862
Rwpos95_82 in95 sp82 3183.098862
Rwpos95_83 in95 sp83 11140.846016
Rwpos95_84 in95 sp84 11140.846016
Rwpos95_85 in95 sp85 3183.098862
Rwpos95_86 in95 sp86 3183.098862
Rwpos95_87 in95 sp87 3183.098862
Rwpos95_88 in95 sp88 3183.098862
Rwpos95_89 in95 sp89 11140.846016
Rwpos95_90 in95 sp90 3183.098862
Rwpos95_91 in95 sp91 11140.846016
Rwpos95_92 in95 sp92 3183.098862
Rwpos95_93 in95 sp93 11140.846016
Rwpos95_94 in95 sp94 11140.846016
Rwpos95_95 in95 sp95 3183.098862
Rwpos95_96 in95 sp96 3183.098862
Rwpos95_97 in95 sp97 11140.846016
Rwpos95_98 in95 sp98 3183.098862
Rwpos95_99 in95 sp99 11140.846016
Rwpos95_100 in95 sp100 3183.098862
Rwpos96_1 in96 sp1 3183.098862
Rwpos96_2 in96 sp2 11140.846016
Rwpos96_3 in96 sp3 11140.846016
Rwpos96_4 in96 sp4 11140.846016
Rwpos96_5 in96 sp5 11140.846016
Rwpos96_6 in96 sp6 3183.098862
Rwpos96_7 in96 sp7 3183.098862
Rwpos96_8 in96 sp8 3183.098862
Rwpos96_9 in96 sp9 11140.846016
Rwpos96_10 in96 sp10 11140.846016
Rwpos96_11 in96 sp11 3183.098862
Rwpos96_12 in96 sp12 3183.098862
Rwpos96_13 in96 sp13 11140.846016
Rwpos96_14 in96 sp14 3183.098862
Rwpos96_15 in96 sp15 11140.846016
Rwpos96_16 in96 sp16 3183.098862
Rwpos96_17 in96 sp17 11140.846016
Rwpos96_18 in96 sp18 11140.846016
Rwpos96_19 in96 sp19 3183.098862
Rwpos96_20 in96 sp20 3183.098862
Rwpos96_21 in96 sp21 3183.098862
Rwpos96_22 in96 sp22 3183.098862
Rwpos96_23 in96 sp23 3183.098862
Rwpos96_24 in96 sp24 3183.098862
Rwpos96_25 in96 sp25 11140.846016
Rwpos96_26 in96 sp26 11140.846016
Rwpos96_27 in96 sp27 11140.846016
Rwpos96_28 in96 sp28 3183.098862
Rwpos96_29 in96 sp29 11140.846016
Rwpos96_30 in96 sp30 3183.098862
Rwpos96_31 in96 sp31 11140.846016
Rwpos96_32 in96 sp32 11140.846016
Rwpos96_33 in96 sp33 3183.098862
Rwpos96_34 in96 sp34 11140.846016
Rwpos96_35 in96 sp35 3183.098862
Rwpos96_36 in96 sp36 3183.098862
Rwpos96_37 in96 sp37 3183.098862
Rwpos96_38 in96 sp38 3183.098862
Rwpos96_39 in96 sp39 3183.098862
Rwpos96_40 in96 sp40 11140.846016
Rwpos96_41 in96 sp41 3183.098862
Rwpos96_42 in96 sp42 3183.098862
Rwpos96_43 in96 sp43 11140.846016
Rwpos96_44 in96 sp44 3183.098862
Rwpos96_45 in96 sp45 3183.098862
Rwpos96_46 in96 sp46 3183.098862
Rwpos96_47 in96 sp47 11140.846016
Rwpos96_48 in96 sp48 3183.098862
Rwpos96_49 in96 sp49 11140.846016
Rwpos96_50 in96 sp50 11140.846016
Rwpos96_51 in96 sp51 3183.098862
Rwpos96_52 in96 sp52 11140.846016
Rwpos96_53 in96 sp53 3183.098862
Rwpos96_54 in96 sp54 3183.098862
Rwpos96_55 in96 sp55 3183.098862
Rwpos96_56 in96 sp56 3183.098862
Rwpos96_57 in96 sp57 3183.098862
Rwpos96_58 in96 sp58 3183.098862
Rwpos96_59 in96 sp59 11140.846016
Rwpos96_60 in96 sp60 3183.098862
Rwpos96_61 in96 sp61 11140.846016
Rwpos96_62 in96 sp62 3183.098862
Rwpos96_63 in96 sp63 11140.846016
Rwpos96_64 in96 sp64 11140.846016
Rwpos96_65 in96 sp65 11140.846016
Rwpos96_66 in96 sp66 3183.098862
Rwpos96_67 in96 sp67 3183.098862
Rwpos96_68 in96 sp68 11140.846016
Rwpos96_69 in96 sp69 11140.846016
Rwpos96_70 in96 sp70 3183.098862
Rwpos96_71 in96 sp71 3183.098862
Rwpos96_72 in96 sp72 3183.098862
Rwpos96_73 in96 sp73 3183.098862
Rwpos96_74 in96 sp74 3183.098862
Rwpos96_75 in96 sp75 11140.846016
Rwpos96_76 in96 sp76 3183.098862
Rwpos96_77 in96 sp77 11140.846016
Rwpos96_78 in96 sp78 3183.098862
Rwpos96_79 in96 sp79 3183.098862
Rwpos96_80 in96 sp80 3183.098862
Rwpos96_81 in96 sp81 11140.846016
Rwpos96_82 in96 sp82 3183.098862
Rwpos96_83 in96 sp83 11140.846016
Rwpos96_84 in96 sp84 3183.098862
Rwpos96_85 in96 sp85 3183.098862
Rwpos96_86 in96 sp86 3183.098862
Rwpos96_87 in96 sp87 3183.098862
Rwpos96_88 in96 sp88 3183.098862
Rwpos96_89 in96 sp89 3183.098862
Rwpos96_90 in96 sp90 3183.098862
Rwpos96_91 in96 sp91 3183.098862
Rwpos96_92 in96 sp92 3183.098862
Rwpos96_93 in96 sp93 11140.846016
Rwpos96_94 in96 sp94 11140.846016
Rwpos96_95 in96 sp95 3183.098862
Rwpos96_96 in96 sp96 11140.846016
Rwpos96_97 in96 sp97 3183.098862
Rwpos96_98 in96 sp98 11140.846016
Rwpos96_99 in96 sp99 11140.846016
Rwpos96_100 in96 sp100 11140.846016
Rwpos97_1 in97 sp1 11140.846016
Rwpos97_2 in97 sp2 3183.098862
Rwpos97_3 in97 sp3 3183.098862
Rwpos97_4 in97 sp4 3183.098862
Rwpos97_5 in97 sp5 11140.846016
Rwpos97_6 in97 sp6 11140.846016
Rwpos97_7 in97 sp7 11140.846016
Rwpos97_8 in97 sp8 3183.098862
Rwpos97_9 in97 sp9 11140.846016
Rwpos97_10 in97 sp10 11140.846016
Rwpos97_11 in97 sp11 3183.098862
Rwpos97_12 in97 sp12 3183.098862
Rwpos97_13 in97 sp13 11140.846016
Rwpos97_14 in97 sp14 3183.098862
Rwpos97_15 in97 sp15 11140.846016
Rwpos97_16 in97 sp16 11140.846016
Rwpos97_17 in97 sp17 11140.846016
Rwpos97_18 in97 sp18 3183.098862
Rwpos97_19 in97 sp19 3183.098862
Rwpos97_20 in97 sp20 11140.846016
Rwpos97_21 in97 sp21 11140.846016
Rwpos97_22 in97 sp22 11140.846016
Rwpos97_23 in97 sp23 3183.098862
Rwpos97_24 in97 sp24 3183.098862
Rwpos97_25 in97 sp25 3183.098862
Rwpos97_26 in97 sp26 11140.846016
Rwpos97_27 in97 sp27 3183.098862
Rwpos97_28 in97 sp28 11140.846016
Rwpos97_29 in97 sp29 3183.098862
Rwpos97_30 in97 sp30 3183.098862
Rwpos97_31 in97 sp31 11140.846016
Rwpos97_32 in97 sp32 11140.846016
Rwpos97_33 in97 sp33 3183.098862
Rwpos97_34 in97 sp34 3183.098862
Rwpos97_35 in97 sp35 3183.098862
Rwpos97_36 in97 sp36 3183.098862
Rwpos97_37 in97 sp37 3183.098862
Rwpos97_38 in97 sp38 11140.846016
Rwpos97_39 in97 sp39 11140.846016
Rwpos97_40 in97 sp40 3183.098862
Rwpos97_41 in97 sp41 11140.846016
Rwpos97_42 in97 sp42 11140.846016
Rwpos97_43 in97 sp43 3183.098862
Rwpos97_44 in97 sp44 3183.098862
Rwpos97_45 in97 sp45 3183.098862
Rwpos97_46 in97 sp46 11140.846016
Rwpos97_47 in97 sp47 11140.846016
Rwpos97_48 in97 sp48 3183.098862
Rwpos97_49 in97 sp49 11140.846016
Rwpos97_50 in97 sp50 3183.098862
Rwpos97_51 in97 sp51 3183.098862
Rwpos97_52 in97 sp52 11140.846016
Rwpos97_53 in97 sp53 11140.846016
Rwpos97_54 in97 sp54 11140.846016
Rwpos97_55 in97 sp55 11140.846016
Rwpos97_56 in97 sp56 3183.098862
Rwpos97_57 in97 sp57 3183.098862
Rwpos97_58 in97 sp58 11140.846016
Rwpos97_59 in97 sp59 3183.098862
Rwpos97_60 in97 sp60 11140.846016
Rwpos97_61 in97 sp61 3183.098862
Rwpos97_62 in97 sp62 11140.846016
Rwpos97_63 in97 sp63 3183.098862
Rwpos97_64 in97 sp64 11140.846016
Rwpos97_65 in97 sp65 3183.098862
Rwpos97_66 in97 sp66 11140.846016
Rwpos97_67 in97 sp67 3183.098862
Rwpos97_68 in97 sp68 11140.846016
Rwpos97_69 in97 sp69 11140.846016
Rwpos97_70 in97 sp70 11140.846016
Rwpos97_71 in97 sp71 11140.846016
Rwpos97_72 in97 sp72 3183.098862
Rwpos97_73 in97 sp73 11140.846016
Rwpos97_74 in97 sp74 3183.098862
Rwpos97_75 in97 sp75 3183.098862
Rwpos97_76 in97 sp76 3183.098862
Rwpos97_77 in97 sp77 3183.098862
Rwpos97_78 in97 sp78 3183.098862
Rwpos97_79 in97 sp79 3183.098862
Rwpos97_80 in97 sp80 11140.846016
Rwpos97_81 in97 sp81 11140.846016
Rwpos97_82 in97 sp82 11140.846016
Rwpos97_83 in97 sp83 3183.098862
Rwpos97_84 in97 sp84 3183.098862
Rwpos97_85 in97 sp85 3183.098862
Rwpos97_86 in97 sp86 3183.098862
Rwpos97_87 in97 sp87 11140.846016
Rwpos97_88 in97 sp88 11140.846016
Rwpos97_89 in97 sp89 3183.098862
Rwpos97_90 in97 sp90 11140.846016
Rwpos97_91 in97 sp91 11140.846016
Rwpos97_92 in97 sp92 11140.846016
Rwpos97_93 in97 sp93 3183.098862
Rwpos97_94 in97 sp94 11140.846016
Rwpos97_95 in97 sp95 3183.098862
Rwpos97_96 in97 sp96 11140.846016
Rwpos97_97 in97 sp97 11140.846016
Rwpos97_98 in97 sp98 11140.846016
Rwpos97_99 in97 sp99 3183.098862
Rwpos97_100 in97 sp100 3183.098862
Rwpos98_1 in98 sp1 11140.846016
Rwpos98_2 in98 sp2 11140.846016
Rwpos98_3 in98 sp3 11140.846016
Rwpos98_4 in98 sp4 3183.098862
Rwpos98_5 in98 sp5 3183.098862
Rwpos98_6 in98 sp6 11140.846016
Rwpos98_7 in98 sp7 3183.098862
Rwpos98_8 in98 sp8 11140.846016
Rwpos98_9 in98 sp9 3183.098862
Rwpos98_10 in98 sp10 3183.098862
Rwpos98_11 in98 sp11 3183.098862
Rwpos98_12 in98 sp12 11140.846016
Rwpos98_13 in98 sp13 11140.846016
Rwpos98_14 in98 sp14 3183.098862
Rwpos98_15 in98 sp15 11140.846016
Rwpos98_16 in98 sp16 3183.098862
Rwpos98_17 in98 sp17 3183.098862
Rwpos98_18 in98 sp18 3183.098862
Rwpos98_19 in98 sp19 3183.098862
Rwpos98_20 in98 sp20 3183.098862
Rwpos98_21 in98 sp21 11140.846016
Rwpos98_22 in98 sp22 3183.098862
Rwpos98_23 in98 sp23 11140.846016
Rwpos98_24 in98 sp24 11140.846016
Rwpos98_25 in98 sp25 11140.846016
Rwpos98_26 in98 sp26 11140.846016
Rwpos98_27 in98 sp27 3183.098862
Rwpos98_28 in98 sp28 11140.846016
Rwpos98_29 in98 sp29 11140.846016
Rwpos98_30 in98 sp30 3183.098862
Rwpos98_31 in98 sp31 3183.098862
Rwpos98_32 in98 sp32 3183.098862
Rwpos98_33 in98 sp33 11140.846016
Rwpos98_34 in98 sp34 3183.098862
Rwpos98_35 in98 sp35 3183.098862
Rwpos98_36 in98 sp36 11140.846016
Rwpos98_37 in98 sp37 11140.846016
Rwpos98_38 in98 sp38 3183.098862
Rwpos98_39 in98 sp39 11140.846016
Rwpos98_40 in98 sp40 3183.098862
Rwpos98_41 in98 sp41 11140.846016
Rwpos98_42 in98 sp42 3183.098862
Rwpos98_43 in98 sp43 3183.098862
Rwpos98_44 in98 sp44 3183.098862
Rwpos98_45 in98 sp45 3183.098862
Rwpos98_46 in98 sp46 3183.098862
Rwpos98_47 in98 sp47 11140.846016
Rwpos98_48 in98 sp48 3183.098862
Rwpos98_49 in98 sp49 3183.098862
Rwpos98_50 in98 sp50 3183.098862
Rwpos98_51 in98 sp51 3183.098862
Rwpos98_52 in98 sp52 11140.846016
Rwpos98_53 in98 sp53 11140.846016
Rwpos98_54 in98 sp54 3183.098862
Rwpos98_55 in98 sp55 3183.098862
Rwpos98_56 in98 sp56 11140.846016
Rwpos98_57 in98 sp57 3183.098862
Rwpos98_58 in98 sp58 11140.846016
Rwpos98_59 in98 sp59 11140.846016
Rwpos98_60 in98 sp60 11140.846016
Rwpos98_61 in98 sp61 3183.098862
Rwpos98_62 in98 sp62 3183.098862
Rwpos98_63 in98 sp63 11140.846016
Rwpos98_64 in98 sp64 3183.098862
Rwpos98_65 in98 sp65 11140.846016
Rwpos98_66 in98 sp66 3183.098862
Rwpos98_67 in98 sp67 11140.846016
Rwpos98_68 in98 sp68 3183.098862
Rwpos98_69 in98 sp69 3183.098862
Rwpos98_70 in98 sp70 3183.098862
Rwpos98_71 in98 sp71 11140.846016
Rwpos98_72 in98 sp72 11140.846016
Rwpos98_73 in98 sp73 3183.098862
Rwpos98_74 in98 sp74 11140.846016
Rwpos98_75 in98 sp75 3183.098862
Rwpos98_76 in98 sp76 11140.846016
Rwpos98_77 in98 sp77 3183.098862
Rwpos98_78 in98 sp78 11140.846016
Rwpos98_79 in98 sp79 3183.098862
Rwpos98_80 in98 sp80 11140.846016
Rwpos98_81 in98 sp81 11140.846016
Rwpos98_82 in98 sp82 3183.098862
Rwpos98_83 in98 sp83 11140.846016
Rwpos98_84 in98 sp84 11140.846016
Rwpos98_85 in98 sp85 11140.846016
Rwpos98_86 in98 sp86 3183.098862
Rwpos98_87 in98 sp87 11140.846016
Rwpos98_88 in98 sp88 11140.846016
Rwpos98_89 in98 sp89 11140.846016
Rwpos98_90 in98 sp90 11140.846016
Rwpos98_91 in98 sp91 11140.846016
Rwpos98_92 in98 sp92 11140.846016
Rwpos98_93 in98 sp93 3183.098862
Rwpos98_94 in98 sp94 11140.846016
Rwpos98_95 in98 sp95 3183.098862
Rwpos98_96 in98 sp96 11140.846016
Rwpos98_97 in98 sp97 11140.846016
Rwpos98_98 in98 sp98 3183.098862
Rwpos98_99 in98 sp99 11140.846016
Rwpos98_100 in98 sp100 3183.098862
Rwpos99_1 in99 sp1 3183.098862
Rwpos99_2 in99 sp2 11140.846016
Rwpos99_3 in99 sp3 11140.846016
Rwpos99_4 in99 sp4 11140.846016
Rwpos99_5 in99 sp5 11140.846016
Rwpos99_6 in99 sp6 11140.846016
Rwpos99_7 in99 sp7 3183.098862
Rwpos99_8 in99 sp8 11140.846016
Rwpos99_9 in99 sp9 3183.098862
Rwpos99_10 in99 sp10 11140.846016
Rwpos99_11 in99 sp11 3183.098862
Rwpos99_12 in99 sp12 11140.846016
Rwpos99_13 in99 sp13 3183.098862
Rwpos99_14 in99 sp14 11140.846016
Rwpos99_15 in99 sp15 3183.098862
Rwpos99_16 in99 sp16 3183.098862
Rwpos99_17 in99 sp17 3183.098862
Rwpos99_18 in99 sp18 3183.098862
Rwpos99_19 in99 sp19 11140.846016
Rwpos99_20 in99 sp20 11140.846016
Rwpos99_21 in99 sp21 3183.098862
Rwpos99_22 in99 sp22 11140.846016
Rwpos99_23 in99 sp23 11140.846016
Rwpos99_24 in99 sp24 11140.846016
Rwpos99_25 in99 sp25 3183.098862
Rwpos99_26 in99 sp26 3183.098862
Rwpos99_27 in99 sp27 11140.846016
Rwpos99_28 in99 sp28 11140.846016
Rwpos99_29 in99 sp29 11140.846016
Rwpos99_30 in99 sp30 11140.846016
Rwpos99_31 in99 sp31 11140.846016
Rwpos99_32 in99 sp32 11140.846016
Rwpos99_33 in99 sp33 11140.846016
Rwpos99_34 in99 sp34 11140.846016
Rwpos99_35 in99 sp35 11140.846016
Rwpos99_36 in99 sp36 3183.098862
Rwpos99_37 in99 sp37 11140.846016
Rwpos99_38 in99 sp38 11140.846016
Rwpos99_39 in99 sp39 3183.098862
Rwpos99_40 in99 sp40 3183.098862
Rwpos99_41 in99 sp41 3183.098862
Rwpos99_42 in99 sp42 11140.846016
Rwpos99_43 in99 sp43 3183.098862
Rwpos99_44 in99 sp44 3183.098862
Rwpos99_45 in99 sp45 3183.098862
Rwpos99_46 in99 sp46 11140.846016
Rwpos99_47 in99 sp47 3183.098862
Rwpos99_48 in99 sp48 3183.098862
Rwpos99_49 in99 sp49 3183.098862
Rwpos99_50 in99 sp50 11140.846016
Rwpos99_51 in99 sp51 3183.098862
Rwpos99_52 in99 sp52 11140.846016
Rwpos99_53 in99 sp53 3183.098862
Rwpos99_54 in99 sp54 11140.846016
Rwpos99_55 in99 sp55 11140.846016
Rwpos99_56 in99 sp56 3183.098862
Rwpos99_57 in99 sp57 11140.846016
Rwpos99_58 in99 sp58 11140.846016
Rwpos99_59 in99 sp59 11140.846016
Rwpos99_60 in99 sp60 11140.846016
Rwpos99_61 in99 sp61 3183.098862
Rwpos99_62 in99 sp62 11140.846016
Rwpos99_63 in99 sp63 11140.846016
Rwpos99_64 in99 sp64 11140.846016
Rwpos99_65 in99 sp65 3183.098862
Rwpos99_66 in99 sp66 11140.846016
Rwpos99_67 in99 sp67 11140.846016
Rwpos99_68 in99 sp68 3183.098862
Rwpos99_69 in99 sp69 11140.846016
Rwpos99_70 in99 sp70 11140.846016
Rwpos99_71 in99 sp71 3183.098862
Rwpos99_72 in99 sp72 11140.846016
Rwpos99_73 in99 sp73 11140.846016
Rwpos99_74 in99 sp74 3183.098862
Rwpos99_75 in99 sp75 3183.098862
Rwpos99_76 in99 sp76 3183.098862
Rwpos99_77 in99 sp77 11140.846016
Rwpos99_78 in99 sp78 3183.098862
Rwpos99_79 in99 sp79 3183.098862
Rwpos99_80 in99 sp80 3183.098862
Rwpos99_81 in99 sp81 3183.098862
Rwpos99_82 in99 sp82 3183.098862
Rwpos99_83 in99 sp83 3183.098862
Rwpos99_84 in99 sp84 3183.098862
Rwpos99_85 in99 sp85 11140.846016
Rwpos99_86 in99 sp86 11140.846016
Rwpos99_87 in99 sp87 3183.098862
Rwpos99_88 in99 sp88 11140.846016
Rwpos99_89 in99 sp89 3183.098862
Rwpos99_90 in99 sp90 11140.846016
Rwpos99_91 in99 sp91 3183.098862
Rwpos99_92 in99 sp92 3183.098862
Rwpos99_93 in99 sp93 11140.846016
Rwpos99_94 in99 sp94 11140.846016
Rwpos99_95 in99 sp95 11140.846016
Rwpos99_96 in99 sp96 3183.098862
Rwpos99_97 in99 sp97 11140.846016
Rwpos99_98 in99 sp98 3183.098862
Rwpos99_99 in99 sp99 11140.846016
Rwpos99_100 in99 sp100 11140.846016
Rwpos100_1 in100 sp1 11140.846016
Rwpos100_2 in100 sp2 11140.846016
Rwpos100_3 in100 sp3 11140.846016
Rwpos100_4 in100 sp4 11140.846016
Rwpos100_5 in100 sp5 11140.846016
Rwpos100_6 in100 sp6 11140.846016
Rwpos100_7 in100 sp7 3183.098862
Rwpos100_8 in100 sp8 11140.846016
Rwpos100_9 in100 sp9 11140.846016
Rwpos100_10 in100 sp10 3183.098862
Rwpos100_11 in100 sp11 3183.098862
Rwpos100_12 in100 sp12 3183.098862
Rwpos100_13 in100 sp13 3183.098862
Rwpos100_14 in100 sp14 11140.846016
Rwpos100_15 in100 sp15 11140.846016
Rwpos100_16 in100 sp16 11140.846016
Rwpos100_17 in100 sp17 3183.098862
Rwpos100_18 in100 sp18 3183.098862
Rwpos100_19 in100 sp19 3183.098862
Rwpos100_20 in100 sp20 3183.098862
Rwpos100_21 in100 sp21 11140.846016
Rwpos100_22 in100 sp22 3183.098862
Rwpos100_23 in100 sp23 3183.098862
Rwpos100_24 in100 sp24 3183.098862
Rwpos100_25 in100 sp25 11140.846016
Rwpos100_26 in100 sp26 11140.846016
Rwpos100_27 in100 sp27 3183.098862
Rwpos100_28 in100 sp28 3183.098862
Rwpos100_29 in100 sp29 3183.098862
Rwpos100_30 in100 sp30 3183.098862
Rwpos100_31 in100 sp31 11140.846016
Rwpos100_32 in100 sp32 3183.098862
Rwpos100_33 in100 sp33 3183.098862
Rwpos100_34 in100 sp34 3183.098862
Rwpos100_35 in100 sp35 3183.098862
Rwpos100_36 in100 sp36 3183.098862
Rwpos100_37 in100 sp37 11140.846016
Rwpos100_38 in100 sp38 3183.098862
Rwpos100_39 in100 sp39 3183.098862
Rwpos100_40 in100 sp40 3183.098862
Rwpos100_41 in100 sp41 3183.098862
Rwpos100_42 in100 sp42 11140.846016
Rwpos100_43 in100 sp43 11140.846016
Rwpos100_44 in100 sp44 3183.098862
Rwpos100_45 in100 sp45 3183.098862
Rwpos100_46 in100 sp46 11140.846016
Rwpos100_47 in100 sp47 11140.846016
Rwpos100_48 in100 sp48 11140.846016
Rwpos100_49 in100 sp49 3183.098862
Rwpos100_50 in100 sp50 3183.098862
Rwpos100_51 in100 sp51 11140.846016
Rwpos100_52 in100 sp52 11140.846016
Rwpos100_53 in100 sp53 3183.098862
Rwpos100_54 in100 sp54 11140.846016
Rwpos100_55 in100 sp55 3183.098862
Rwpos100_56 in100 sp56 11140.846016
Rwpos100_57 in100 sp57 3183.098862
Rwpos100_58 in100 sp58 11140.846016
Rwpos100_59 in100 sp59 11140.846016
Rwpos100_60 in100 sp60 3183.098862
Rwpos100_61 in100 sp61 3183.098862
Rwpos100_62 in100 sp62 3183.098862
Rwpos100_63 in100 sp63 11140.846016
Rwpos100_64 in100 sp64 11140.846016
Rwpos100_65 in100 sp65 3183.098862
Rwpos100_66 in100 sp66 11140.846016
Rwpos100_67 in100 sp67 3183.098862
Rwpos100_68 in100 sp68 11140.846016
Rwpos100_69 in100 sp69 11140.846016
Rwpos100_70 in100 sp70 11140.846016
Rwpos100_71 in100 sp71 3183.098862
Rwpos100_72 in100 sp72 3183.098862
Rwpos100_73 in100 sp73 3183.098862
Rwpos100_74 in100 sp74 3183.098862
Rwpos100_75 in100 sp75 3183.098862
Rwpos100_76 in100 sp76 3183.098862
Rwpos100_77 in100 sp77 3183.098862
Rwpos100_78 in100 sp78 3183.098862
Rwpos100_79 in100 sp79 11140.846016
Rwpos100_80 in100 sp80 11140.846016
Rwpos100_81 in100 sp81 11140.846016
Rwpos100_82 in100 sp82 3183.098862
Rwpos100_83 in100 sp83 3183.098862
Rwpos100_84 in100 sp84 3183.098862
Rwpos100_85 in100 sp85 3183.098862
Rwpos100_86 in100 sp86 11140.846016
Rwpos100_87 in100 sp87 3183.098862
Rwpos100_88 in100 sp88 11140.846016
Rwpos100_89 in100 sp89 11140.846016
Rwpos100_90 in100 sp90 11140.846016
Rwpos100_91 in100 sp91 11140.846016
Rwpos100_92 in100 sp92 3183.098862
Rwpos100_93 in100 sp93 11140.846016
Rwpos100_94 in100 sp94 3183.098862
Rwpos100_95 in100 sp95 3183.098862
Rwpos100_96 in100 sp96 11140.846016
Rwpos100_97 in100 sp97 3183.098862
Rwpos100_98 in100 sp98 3183.098862
Rwpos100_99 in100 sp99 11140.846016
Rwpos100_100 in100 sp100 11140.846016
Rwpos101_1 in101 sp1 11140.846016
Rwpos101_2 in101 sp2 3183.098862
Rwpos101_3 in101 sp3 3183.098862
Rwpos101_4 in101 sp4 11140.846016
Rwpos101_5 in101 sp5 3183.098862
Rwpos101_6 in101 sp6 11140.846016
Rwpos101_7 in101 sp7 11140.846016
Rwpos101_8 in101 sp8 3183.098862
Rwpos101_9 in101 sp9 11140.846016
Rwpos101_10 in101 sp10 3183.098862
Rwpos101_11 in101 sp11 11140.846016
Rwpos101_12 in101 sp12 11140.846016
Rwpos101_13 in101 sp13 11140.846016
Rwpos101_14 in101 sp14 3183.098862
Rwpos101_15 in101 sp15 11140.846016
Rwpos101_16 in101 sp16 3183.098862
Rwpos101_17 in101 sp17 3183.098862
Rwpos101_18 in101 sp18 3183.098862
Rwpos101_19 in101 sp19 3183.098862
Rwpos101_20 in101 sp20 3183.098862
Rwpos101_21 in101 sp21 3183.098862
Rwpos101_22 in101 sp22 3183.098862
Rwpos101_23 in101 sp23 11140.846016
Rwpos101_24 in101 sp24 3183.098862
Rwpos101_25 in101 sp25 11140.846016
Rwpos101_26 in101 sp26 3183.098862
Rwpos101_27 in101 sp27 3183.098862
Rwpos101_28 in101 sp28 11140.846016
Rwpos101_29 in101 sp29 3183.098862
Rwpos101_30 in101 sp30 3183.098862
Rwpos101_31 in101 sp31 11140.846016
Rwpos101_32 in101 sp32 3183.098862
Rwpos101_33 in101 sp33 11140.846016
Rwpos101_34 in101 sp34 11140.846016
Rwpos101_35 in101 sp35 3183.098862
Rwpos101_36 in101 sp36 3183.098862
Rwpos101_37 in101 sp37 3183.098862
Rwpos101_38 in101 sp38 11140.846016
Rwpos101_39 in101 sp39 3183.098862
Rwpos101_40 in101 sp40 3183.098862
Rwpos101_41 in101 sp41 11140.846016
Rwpos101_42 in101 sp42 3183.098862
Rwpos101_43 in101 sp43 3183.098862
Rwpos101_44 in101 sp44 3183.098862
Rwpos101_45 in101 sp45 11140.846016
Rwpos101_46 in101 sp46 3183.098862
Rwpos101_47 in101 sp47 3183.098862
Rwpos101_48 in101 sp48 3183.098862
Rwpos101_49 in101 sp49 3183.098862
Rwpos101_50 in101 sp50 11140.846016
Rwpos101_51 in101 sp51 3183.098862
Rwpos101_52 in101 sp52 3183.098862
Rwpos101_53 in101 sp53 11140.846016
Rwpos101_54 in101 sp54 3183.098862
Rwpos101_55 in101 sp55 3183.098862
Rwpos101_56 in101 sp56 11140.846016
Rwpos101_57 in101 sp57 11140.846016
Rwpos101_58 in101 sp58 3183.098862
Rwpos101_59 in101 sp59 3183.098862
Rwpos101_60 in101 sp60 11140.846016
Rwpos101_61 in101 sp61 11140.846016
Rwpos101_62 in101 sp62 3183.098862
Rwpos101_63 in101 sp63 11140.846016
Rwpos101_64 in101 sp64 3183.098862
Rwpos101_65 in101 sp65 11140.846016
Rwpos101_66 in101 sp66 11140.846016
Rwpos101_67 in101 sp67 3183.098862
Rwpos101_68 in101 sp68 3183.098862
Rwpos101_69 in101 sp69 11140.846016
Rwpos101_70 in101 sp70 3183.098862
Rwpos101_71 in101 sp71 3183.098862
Rwpos101_72 in101 sp72 11140.846016
Rwpos101_73 in101 sp73 11140.846016
Rwpos101_74 in101 sp74 3183.098862
Rwpos101_75 in101 sp75 3183.098862
Rwpos101_76 in101 sp76 3183.098862
Rwpos101_77 in101 sp77 11140.846016
Rwpos101_78 in101 sp78 11140.846016
Rwpos101_79 in101 sp79 11140.846016
Rwpos101_80 in101 sp80 3183.098862
Rwpos101_81 in101 sp81 11140.846016
Rwpos101_82 in101 sp82 11140.846016
Rwpos101_83 in101 sp83 3183.098862
Rwpos101_84 in101 sp84 3183.098862
Rwpos101_85 in101 sp85 3183.098862
Rwpos101_86 in101 sp86 3183.098862
Rwpos101_87 in101 sp87 3183.098862
Rwpos101_88 in101 sp88 3183.098862
Rwpos101_89 in101 sp89 3183.098862
Rwpos101_90 in101 sp90 11140.846016
Rwpos101_91 in101 sp91 3183.098862
Rwpos101_92 in101 sp92 11140.846016
Rwpos101_93 in101 sp93 11140.846016
Rwpos101_94 in101 sp94 3183.098862
Rwpos101_95 in101 sp95 11140.846016
Rwpos101_96 in101 sp96 3183.098862
Rwpos101_97 in101 sp97 11140.846016
Rwpos101_98 in101 sp98 11140.846016
Rwpos101_99 in101 sp99 3183.098862
Rwpos101_100 in101 sp100 11140.846016
Rwpos102_1 in102 sp1 3183.098862
Rwpos102_2 in102 sp2 3183.098862
Rwpos102_3 in102 sp3 11140.846016
Rwpos102_4 in102 sp4 11140.846016
Rwpos102_5 in102 sp5 11140.846016
Rwpos102_6 in102 sp6 3183.098862
Rwpos102_7 in102 sp7 3183.098862
Rwpos102_8 in102 sp8 3183.098862
Rwpos102_9 in102 sp9 11140.846016
Rwpos102_10 in102 sp10 11140.846016
Rwpos102_11 in102 sp11 11140.846016
Rwpos102_12 in102 sp12 3183.098862
Rwpos102_13 in102 sp13 3183.098862
Rwpos102_14 in102 sp14 11140.846016
Rwpos102_15 in102 sp15 3183.098862
Rwpos102_16 in102 sp16 11140.846016
Rwpos102_17 in102 sp17 11140.846016
Rwpos102_18 in102 sp18 11140.846016
Rwpos102_19 in102 sp19 11140.846016
Rwpos102_20 in102 sp20 11140.846016
Rwpos102_21 in102 sp21 11140.846016
Rwpos102_22 in102 sp22 11140.846016
Rwpos102_23 in102 sp23 3183.098862
Rwpos102_24 in102 sp24 3183.098862
Rwpos102_25 in102 sp25 3183.098862
Rwpos102_26 in102 sp26 3183.098862
Rwpos102_27 in102 sp27 3183.098862
Rwpos102_28 in102 sp28 3183.098862
Rwpos102_29 in102 sp29 3183.098862
Rwpos102_30 in102 sp30 3183.098862
Rwpos102_31 in102 sp31 3183.098862
Rwpos102_32 in102 sp32 3183.098862
Rwpos102_33 in102 sp33 3183.098862
Rwpos102_34 in102 sp34 3183.098862
Rwpos102_35 in102 sp35 11140.846016
Rwpos102_36 in102 sp36 3183.098862
Rwpos102_37 in102 sp37 11140.846016
Rwpos102_38 in102 sp38 3183.098862
Rwpos102_39 in102 sp39 11140.846016
Rwpos102_40 in102 sp40 3183.098862
Rwpos102_41 in102 sp41 11140.846016
Rwpos102_42 in102 sp42 11140.846016
Rwpos102_43 in102 sp43 3183.098862
Rwpos102_44 in102 sp44 11140.846016
Rwpos102_45 in102 sp45 3183.098862
Rwpos102_46 in102 sp46 11140.846016
Rwpos102_47 in102 sp47 3183.098862
Rwpos102_48 in102 sp48 11140.846016
Rwpos102_49 in102 sp49 11140.846016
Rwpos102_50 in102 sp50 11140.846016
Rwpos102_51 in102 sp51 3183.098862
Rwpos102_52 in102 sp52 11140.846016
Rwpos102_53 in102 sp53 11140.846016
Rwpos102_54 in102 sp54 3183.098862
Rwpos102_55 in102 sp55 11140.846016
Rwpos102_56 in102 sp56 3183.098862
Rwpos102_57 in102 sp57 3183.098862
Rwpos102_58 in102 sp58 11140.846016
Rwpos102_59 in102 sp59 3183.098862
Rwpos102_60 in102 sp60 11140.846016
Rwpos102_61 in102 sp61 11140.846016
Rwpos102_62 in102 sp62 11140.846016
Rwpos102_63 in102 sp63 3183.098862
Rwpos102_64 in102 sp64 3183.098862
Rwpos102_65 in102 sp65 3183.098862
Rwpos102_66 in102 sp66 11140.846016
Rwpos102_67 in102 sp67 3183.098862
Rwpos102_68 in102 sp68 3183.098862
Rwpos102_69 in102 sp69 11140.846016
Rwpos102_70 in102 sp70 11140.846016
Rwpos102_71 in102 sp71 11140.846016
Rwpos102_72 in102 sp72 11140.846016
Rwpos102_73 in102 sp73 11140.846016
Rwpos102_74 in102 sp74 3183.098862
Rwpos102_75 in102 sp75 3183.098862
Rwpos102_76 in102 sp76 11140.846016
Rwpos102_77 in102 sp77 3183.098862
Rwpos102_78 in102 sp78 11140.846016
Rwpos102_79 in102 sp79 3183.098862
Rwpos102_80 in102 sp80 3183.098862
Rwpos102_81 in102 sp81 3183.098862
Rwpos102_82 in102 sp82 3183.098862
Rwpos102_83 in102 sp83 3183.098862
Rwpos102_84 in102 sp84 3183.098862
Rwpos102_85 in102 sp85 3183.098862
Rwpos102_86 in102 sp86 3183.098862
Rwpos102_87 in102 sp87 11140.846016
Rwpos102_88 in102 sp88 11140.846016
Rwpos102_89 in102 sp89 11140.846016
Rwpos102_90 in102 sp90 11140.846016
Rwpos102_91 in102 sp91 3183.098862
Rwpos102_92 in102 sp92 11140.846016
Rwpos102_93 in102 sp93 11140.846016
Rwpos102_94 in102 sp94 3183.098862
Rwpos102_95 in102 sp95 3183.098862
Rwpos102_96 in102 sp96 3183.098862
Rwpos102_97 in102 sp97 3183.098862
Rwpos102_98 in102 sp98 11140.846016
Rwpos102_99 in102 sp99 11140.846016
Rwpos102_100 in102 sp100 3183.098862
Rwpos103_1 in103 sp1 11140.846016
Rwpos103_2 in103 sp2 3183.098862
Rwpos103_3 in103 sp3 11140.846016
Rwpos103_4 in103 sp4 11140.846016
Rwpos103_5 in103 sp5 11140.846016
Rwpos103_6 in103 sp6 11140.846016
Rwpos103_7 in103 sp7 3183.098862
Rwpos103_8 in103 sp8 11140.846016
Rwpos103_9 in103 sp9 3183.098862
Rwpos103_10 in103 sp10 11140.846016
Rwpos103_11 in103 sp11 3183.098862
Rwpos103_12 in103 sp12 3183.098862
Rwpos103_13 in103 sp13 11140.846016
Rwpos103_14 in103 sp14 3183.098862
Rwpos103_15 in103 sp15 11140.846016
Rwpos103_16 in103 sp16 11140.846016
Rwpos103_17 in103 sp17 11140.846016
Rwpos103_18 in103 sp18 3183.098862
Rwpos103_19 in103 sp19 11140.846016
Rwpos103_20 in103 sp20 11140.846016
Rwpos103_21 in103 sp21 3183.098862
Rwpos103_22 in103 sp22 11140.846016
Rwpos103_23 in103 sp23 3183.098862
Rwpos103_24 in103 sp24 11140.846016
Rwpos103_25 in103 sp25 11140.846016
Rwpos103_26 in103 sp26 3183.098862
Rwpos103_27 in103 sp27 11140.846016
Rwpos103_28 in103 sp28 3183.098862
Rwpos103_29 in103 sp29 11140.846016
Rwpos103_30 in103 sp30 3183.098862
Rwpos103_31 in103 sp31 3183.098862
Rwpos103_32 in103 sp32 11140.846016
Rwpos103_33 in103 sp33 3183.098862
Rwpos103_34 in103 sp34 11140.846016
Rwpos103_35 in103 sp35 11140.846016
Rwpos103_36 in103 sp36 3183.098862
Rwpos103_37 in103 sp37 3183.098862
Rwpos103_38 in103 sp38 11140.846016
Rwpos103_39 in103 sp39 11140.846016
Rwpos103_40 in103 sp40 11140.846016
Rwpos103_41 in103 sp41 11140.846016
Rwpos103_42 in103 sp42 3183.098862
Rwpos103_43 in103 sp43 11140.846016
Rwpos103_44 in103 sp44 3183.098862
Rwpos103_45 in103 sp45 3183.098862
Rwpos103_46 in103 sp46 3183.098862
Rwpos103_47 in103 sp47 11140.846016
Rwpos103_48 in103 sp48 3183.098862
Rwpos103_49 in103 sp49 11140.846016
Rwpos103_50 in103 sp50 3183.098862
Rwpos103_51 in103 sp51 11140.846016
Rwpos103_52 in103 sp52 11140.846016
Rwpos103_53 in103 sp53 3183.098862
Rwpos103_54 in103 sp54 11140.846016
Rwpos103_55 in103 sp55 3183.098862
Rwpos103_56 in103 sp56 11140.846016
Rwpos103_57 in103 sp57 3183.098862
Rwpos103_58 in103 sp58 11140.846016
Rwpos103_59 in103 sp59 3183.098862
Rwpos103_60 in103 sp60 11140.846016
Rwpos103_61 in103 sp61 3183.098862
Rwpos103_62 in103 sp62 11140.846016
Rwpos103_63 in103 sp63 11140.846016
Rwpos103_64 in103 sp64 11140.846016
Rwpos103_65 in103 sp65 11140.846016
Rwpos103_66 in103 sp66 3183.098862
Rwpos103_67 in103 sp67 3183.098862
Rwpos103_68 in103 sp68 11140.846016
Rwpos103_69 in103 sp69 3183.098862
Rwpos103_70 in103 sp70 11140.846016
Rwpos103_71 in103 sp71 3183.098862
Rwpos103_72 in103 sp72 3183.098862
Rwpos103_73 in103 sp73 3183.098862
Rwpos103_74 in103 sp74 11140.846016
Rwpos103_75 in103 sp75 11140.846016
Rwpos103_76 in103 sp76 11140.846016
Rwpos103_77 in103 sp77 3183.098862
Rwpos103_78 in103 sp78 11140.846016
Rwpos103_79 in103 sp79 3183.098862
Rwpos103_80 in103 sp80 11140.846016
Rwpos103_81 in103 sp81 11140.846016
Rwpos103_82 in103 sp82 3183.098862
Rwpos103_83 in103 sp83 11140.846016
Rwpos103_84 in103 sp84 3183.098862
Rwpos103_85 in103 sp85 11140.846016
Rwpos103_86 in103 sp86 11140.846016
Rwpos103_87 in103 sp87 11140.846016
Rwpos103_88 in103 sp88 3183.098862
Rwpos103_89 in103 sp89 3183.098862
Rwpos103_90 in103 sp90 3183.098862
Rwpos103_91 in103 sp91 11140.846016
Rwpos103_92 in103 sp92 11140.846016
Rwpos103_93 in103 sp93 11140.846016
Rwpos103_94 in103 sp94 11140.846016
Rwpos103_95 in103 sp95 3183.098862
Rwpos103_96 in103 sp96 11140.846016
Rwpos103_97 in103 sp97 11140.846016
Rwpos103_98 in103 sp98 11140.846016
Rwpos103_99 in103 sp99 3183.098862
Rwpos103_100 in103 sp100 3183.098862
Rwpos104_1 in104 sp1 11140.846016
Rwpos104_2 in104 sp2 11140.846016
Rwpos104_3 in104 sp3 3183.098862
Rwpos104_4 in104 sp4 3183.098862
Rwpos104_5 in104 sp5 11140.846016
Rwpos104_6 in104 sp6 11140.846016
Rwpos104_7 in104 sp7 11140.846016
Rwpos104_8 in104 sp8 3183.098862
Rwpos104_9 in104 sp9 3183.098862
Rwpos104_10 in104 sp10 3183.098862
Rwpos104_11 in104 sp11 11140.846016
Rwpos104_12 in104 sp12 3183.098862
Rwpos104_13 in104 sp13 11140.846016
Rwpos104_14 in104 sp14 3183.098862
Rwpos104_15 in104 sp15 11140.846016
Rwpos104_16 in104 sp16 11140.846016
Rwpos104_17 in104 sp17 11140.846016
Rwpos104_18 in104 sp18 11140.846016
Rwpos104_19 in104 sp19 3183.098862
Rwpos104_20 in104 sp20 11140.846016
Rwpos104_21 in104 sp21 11140.846016
Rwpos104_22 in104 sp22 11140.846016
Rwpos104_23 in104 sp23 3183.098862
Rwpos104_24 in104 sp24 11140.846016
Rwpos104_25 in104 sp25 11140.846016
Rwpos104_26 in104 sp26 3183.098862
Rwpos104_27 in104 sp27 3183.098862
Rwpos104_28 in104 sp28 3183.098862
Rwpos104_29 in104 sp29 3183.098862
Rwpos104_30 in104 sp30 11140.846016
Rwpos104_31 in104 sp31 11140.846016
Rwpos104_32 in104 sp32 11140.846016
Rwpos104_33 in104 sp33 11140.846016
Rwpos104_34 in104 sp34 11140.846016
Rwpos104_35 in104 sp35 11140.846016
Rwpos104_36 in104 sp36 11140.846016
Rwpos104_37 in104 sp37 3183.098862
Rwpos104_38 in104 sp38 11140.846016
Rwpos104_39 in104 sp39 11140.846016
Rwpos104_40 in104 sp40 11140.846016
Rwpos104_41 in104 sp41 3183.098862
Rwpos104_42 in104 sp42 11140.846016
Rwpos104_43 in104 sp43 3183.098862
Rwpos104_44 in104 sp44 3183.098862
Rwpos104_45 in104 sp45 11140.846016
Rwpos104_46 in104 sp46 3183.098862
Rwpos104_47 in104 sp47 11140.846016
Rwpos104_48 in104 sp48 3183.098862
Rwpos104_49 in104 sp49 11140.846016
Rwpos104_50 in104 sp50 11140.846016
Rwpos104_51 in104 sp51 3183.098862
Rwpos104_52 in104 sp52 3183.098862
Rwpos104_53 in104 sp53 11140.846016
Rwpos104_54 in104 sp54 11140.846016
Rwpos104_55 in104 sp55 11140.846016
Rwpos104_56 in104 sp56 3183.098862
Rwpos104_57 in104 sp57 3183.098862
Rwpos104_58 in104 sp58 11140.846016
Rwpos104_59 in104 sp59 11140.846016
Rwpos104_60 in104 sp60 3183.098862
Rwpos104_61 in104 sp61 11140.846016
Rwpos104_62 in104 sp62 3183.098862
Rwpos104_63 in104 sp63 3183.098862
Rwpos104_64 in104 sp64 3183.098862
Rwpos104_65 in104 sp65 11140.846016
Rwpos104_66 in104 sp66 11140.846016
Rwpos104_67 in104 sp67 11140.846016
Rwpos104_68 in104 sp68 3183.098862
Rwpos104_69 in104 sp69 11140.846016
Rwpos104_70 in104 sp70 3183.098862
Rwpos104_71 in104 sp71 11140.846016
Rwpos104_72 in104 sp72 3183.098862
Rwpos104_73 in104 sp73 11140.846016
Rwpos104_74 in104 sp74 11140.846016
Rwpos104_75 in104 sp75 3183.098862
Rwpos104_76 in104 sp76 3183.098862
Rwpos104_77 in104 sp77 11140.846016
Rwpos104_78 in104 sp78 3183.098862
Rwpos104_79 in104 sp79 11140.846016
Rwpos104_80 in104 sp80 3183.098862
Rwpos104_81 in104 sp81 3183.098862
Rwpos104_82 in104 sp82 11140.846016
Rwpos104_83 in104 sp83 3183.098862
Rwpos104_84 in104 sp84 11140.846016
Rwpos104_85 in104 sp85 11140.846016
Rwpos104_86 in104 sp86 3183.098862
Rwpos104_87 in104 sp87 3183.098862
Rwpos104_88 in104 sp88 11140.846016
Rwpos104_89 in104 sp89 3183.098862
Rwpos104_90 in104 sp90 11140.846016
Rwpos104_91 in104 sp91 11140.846016
Rwpos104_92 in104 sp92 3183.098862
Rwpos104_93 in104 sp93 11140.846016
Rwpos104_94 in104 sp94 3183.098862
Rwpos104_95 in104 sp95 3183.098862
Rwpos104_96 in104 sp96 11140.846016
Rwpos104_97 in104 sp97 11140.846016
Rwpos104_98 in104 sp98 3183.098862
Rwpos104_99 in104 sp99 3183.098862
Rwpos104_100 in104 sp100 3183.098862
Rwpos105_1 in105 sp1 11140.846016
Rwpos105_2 in105 sp2 3183.098862
Rwpos105_3 in105 sp3 3183.098862
Rwpos105_4 in105 sp4 11140.846016
Rwpos105_5 in105 sp5 3183.098862
Rwpos105_6 in105 sp6 11140.846016
Rwpos105_7 in105 sp7 3183.098862
Rwpos105_8 in105 sp8 11140.846016
Rwpos105_9 in105 sp9 11140.846016
Rwpos105_10 in105 sp10 3183.098862
Rwpos105_11 in105 sp11 11140.846016
Rwpos105_12 in105 sp12 3183.098862
Rwpos105_13 in105 sp13 3183.098862
Rwpos105_14 in105 sp14 3183.098862
Rwpos105_15 in105 sp15 3183.098862
Rwpos105_16 in105 sp16 11140.846016
Rwpos105_17 in105 sp17 11140.846016
Rwpos105_18 in105 sp18 3183.098862
Rwpos105_19 in105 sp19 3183.098862
Rwpos105_20 in105 sp20 11140.846016
Rwpos105_21 in105 sp21 11140.846016
Rwpos105_22 in105 sp22 11140.846016
Rwpos105_23 in105 sp23 11140.846016
Rwpos105_24 in105 sp24 11140.846016
Rwpos105_25 in105 sp25 11140.846016
Rwpos105_26 in105 sp26 3183.098862
Rwpos105_27 in105 sp27 11140.846016
Rwpos105_28 in105 sp28 11140.846016
Rwpos105_29 in105 sp29 3183.098862
Rwpos105_30 in105 sp30 3183.098862
Rwpos105_31 in105 sp31 3183.098862
Rwpos105_32 in105 sp32 11140.846016
Rwpos105_33 in105 sp33 11140.846016
Rwpos105_34 in105 sp34 11140.846016
Rwpos105_35 in105 sp35 3183.098862
Rwpos105_36 in105 sp36 11140.846016
Rwpos105_37 in105 sp37 11140.846016
Rwpos105_38 in105 sp38 3183.098862
Rwpos105_39 in105 sp39 11140.846016
Rwpos105_40 in105 sp40 3183.098862
Rwpos105_41 in105 sp41 11140.846016
Rwpos105_42 in105 sp42 3183.098862
Rwpos105_43 in105 sp43 11140.846016
Rwpos105_44 in105 sp44 3183.098862
Rwpos105_45 in105 sp45 11140.846016
Rwpos105_46 in105 sp46 3183.098862
Rwpos105_47 in105 sp47 11140.846016
Rwpos105_48 in105 sp48 3183.098862
Rwpos105_49 in105 sp49 11140.846016
Rwpos105_50 in105 sp50 3183.098862
Rwpos105_51 in105 sp51 3183.098862
Rwpos105_52 in105 sp52 3183.098862
Rwpos105_53 in105 sp53 11140.846016
Rwpos105_54 in105 sp54 11140.846016
Rwpos105_55 in105 sp55 3183.098862
Rwpos105_56 in105 sp56 3183.098862
Rwpos105_57 in105 sp57 3183.098862
Rwpos105_58 in105 sp58 3183.098862
Rwpos105_59 in105 sp59 3183.098862
Rwpos105_60 in105 sp60 3183.098862
Rwpos105_61 in105 sp61 3183.098862
Rwpos105_62 in105 sp62 11140.846016
Rwpos105_63 in105 sp63 3183.098862
Rwpos105_64 in105 sp64 11140.846016
Rwpos105_65 in105 sp65 11140.846016
Rwpos105_66 in105 sp66 11140.846016
Rwpos105_67 in105 sp67 3183.098862
Rwpos105_68 in105 sp68 11140.846016
Rwpos105_69 in105 sp69 3183.098862
Rwpos105_70 in105 sp70 11140.846016
Rwpos105_71 in105 sp71 11140.846016
Rwpos105_72 in105 sp72 11140.846016
Rwpos105_73 in105 sp73 3183.098862
Rwpos105_74 in105 sp74 3183.098862
Rwpos105_75 in105 sp75 3183.098862
Rwpos105_76 in105 sp76 3183.098862
Rwpos105_77 in105 sp77 11140.846016
Rwpos105_78 in105 sp78 3183.098862
Rwpos105_79 in105 sp79 3183.098862
Rwpos105_80 in105 sp80 11140.846016
Rwpos105_81 in105 sp81 11140.846016
Rwpos105_82 in105 sp82 11140.846016
Rwpos105_83 in105 sp83 3183.098862
Rwpos105_84 in105 sp84 3183.098862
Rwpos105_85 in105 sp85 3183.098862
Rwpos105_86 in105 sp86 3183.098862
Rwpos105_87 in105 sp87 11140.846016
Rwpos105_88 in105 sp88 3183.098862
Rwpos105_89 in105 sp89 3183.098862
Rwpos105_90 in105 sp90 3183.098862
Rwpos105_91 in105 sp91 11140.846016
Rwpos105_92 in105 sp92 11140.846016
Rwpos105_93 in105 sp93 11140.846016
Rwpos105_94 in105 sp94 3183.098862
Rwpos105_95 in105 sp95 11140.846016
Rwpos105_96 in105 sp96 3183.098862
Rwpos105_97 in105 sp97 11140.846016
Rwpos105_98 in105 sp98 11140.846016
Rwpos105_99 in105 sp99 11140.846016
Rwpos105_100 in105 sp100 11140.846016
Rwpos106_1 in106 sp1 3183.098862
Rwpos106_2 in106 sp2 11140.846016
Rwpos106_3 in106 sp3 3183.098862
Rwpos106_4 in106 sp4 3183.098862
Rwpos106_5 in106 sp5 11140.846016
Rwpos106_6 in106 sp6 3183.098862
Rwpos106_7 in106 sp7 3183.098862
Rwpos106_8 in106 sp8 3183.098862
Rwpos106_9 in106 sp9 11140.846016
Rwpos106_10 in106 sp10 11140.846016
Rwpos106_11 in106 sp11 3183.098862
Rwpos106_12 in106 sp12 3183.098862
Rwpos106_13 in106 sp13 11140.846016
Rwpos106_14 in106 sp14 11140.846016
Rwpos106_15 in106 sp15 3183.098862
Rwpos106_16 in106 sp16 3183.098862
Rwpos106_17 in106 sp17 3183.098862
Rwpos106_18 in106 sp18 11140.846016
Rwpos106_19 in106 sp19 11140.846016
Rwpos106_20 in106 sp20 11140.846016
Rwpos106_21 in106 sp21 11140.846016
Rwpos106_22 in106 sp22 3183.098862
Rwpos106_23 in106 sp23 3183.098862
Rwpos106_24 in106 sp24 3183.098862
Rwpos106_25 in106 sp25 11140.846016
Rwpos106_26 in106 sp26 11140.846016
Rwpos106_27 in106 sp27 11140.846016
Rwpos106_28 in106 sp28 3183.098862
Rwpos106_29 in106 sp29 3183.098862
Rwpos106_30 in106 sp30 11140.846016
Rwpos106_31 in106 sp31 3183.098862
Rwpos106_32 in106 sp32 11140.846016
Rwpos106_33 in106 sp33 11140.846016
Rwpos106_34 in106 sp34 3183.098862
Rwpos106_35 in106 sp35 3183.098862
Rwpos106_36 in106 sp36 3183.098862
Rwpos106_37 in106 sp37 11140.846016
Rwpos106_38 in106 sp38 3183.098862
Rwpos106_39 in106 sp39 3183.098862
Rwpos106_40 in106 sp40 3183.098862
Rwpos106_41 in106 sp41 11140.846016
Rwpos106_42 in106 sp42 11140.846016
Rwpos106_43 in106 sp43 11140.846016
Rwpos106_44 in106 sp44 3183.098862
Rwpos106_45 in106 sp45 11140.846016
Rwpos106_46 in106 sp46 11140.846016
Rwpos106_47 in106 sp47 3183.098862
Rwpos106_48 in106 sp48 11140.846016
Rwpos106_49 in106 sp49 3183.098862
Rwpos106_50 in106 sp50 11140.846016
Rwpos106_51 in106 sp51 11140.846016
Rwpos106_52 in106 sp52 3183.098862
Rwpos106_53 in106 sp53 3183.098862
Rwpos106_54 in106 sp54 3183.098862
Rwpos106_55 in106 sp55 3183.098862
Rwpos106_56 in106 sp56 3183.098862
Rwpos106_57 in106 sp57 11140.846016
Rwpos106_58 in106 sp58 11140.846016
Rwpos106_59 in106 sp59 11140.846016
Rwpos106_60 in106 sp60 3183.098862
Rwpos106_61 in106 sp61 3183.098862
Rwpos106_62 in106 sp62 11140.846016
Rwpos106_63 in106 sp63 3183.098862
Rwpos106_64 in106 sp64 3183.098862
Rwpos106_65 in106 sp65 11140.846016
Rwpos106_66 in106 sp66 3183.098862
Rwpos106_67 in106 sp67 11140.846016
Rwpos106_68 in106 sp68 3183.098862
Rwpos106_69 in106 sp69 3183.098862
Rwpos106_70 in106 sp70 11140.846016
Rwpos106_71 in106 sp71 3183.098862
Rwpos106_72 in106 sp72 11140.846016
Rwpos106_73 in106 sp73 11140.846016
Rwpos106_74 in106 sp74 3183.098862
Rwpos106_75 in106 sp75 3183.098862
Rwpos106_76 in106 sp76 3183.098862
Rwpos106_77 in106 sp77 11140.846016
Rwpos106_78 in106 sp78 11140.846016
Rwpos106_79 in106 sp79 3183.098862
Rwpos106_80 in106 sp80 11140.846016
Rwpos106_81 in106 sp81 11140.846016
Rwpos106_82 in106 sp82 3183.098862
Rwpos106_83 in106 sp83 11140.846016
Rwpos106_84 in106 sp84 3183.098862
Rwpos106_85 in106 sp85 11140.846016
Rwpos106_86 in106 sp86 3183.098862
Rwpos106_87 in106 sp87 3183.098862
Rwpos106_88 in106 sp88 3183.098862
Rwpos106_89 in106 sp89 11140.846016
Rwpos106_90 in106 sp90 11140.846016
Rwpos106_91 in106 sp91 11140.846016
Rwpos106_92 in106 sp92 3183.098862
Rwpos106_93 in106 sp93 3183.098862
Rwpos106_94 in106 sp94 11140.846016
Rwpos106_95 in106 sp95 11140.846016
Rwpos106_96 in106 sp96 3183.098862
Rwpos106_97 in106 sp97 3183.098862
Rwpos106_98 in106 sp98 3183.098862
Rwpos106_99 in106 sp99 11140.846016
Rwpos106_100 in106 sp100 11140.846016
Rwpos107_1 in107 sp1 3183.098862
Rwpos107_2 in107 sp2 11140.846016
Rwpos107_3 in107 sp3 3183.098862
Rwpos107_4 in107 sp4 3183.098862
Rwpos107_5 in107 sp5 11140.846016
Rwpos107_6 in107 sp6 3183.098862
Rwpos107_7 in107 sp7 3183.098862
Rwpos107_8 in107 sp8 3183.098862
Rwpos107_9 in107 sp9 3183.098862
Rwpos107_10 in107 sp10 11140.846016
Rwpos107_11 in107 sp11 11140.846016
Rwpos107_12 in107 sp12 3183.098862
Rwpos107_13 in107 sp13 3183.098862
Rwpos107_14 in107 sp14 3183.098862
Rwpos107_15 in107 sp15 3183.098862
Rwpos107_16 in107 sp16 3183.098862
Rwpos107_17 in107 sp17 11140.846016
Rwpos107_18 in107 sp18 3183.098862
Rwpos107_19 in107 sp19 3183.098862
Rwpos107_20 in107 sp20 11140.846016
Rwpos107_21 in107 sp21 11140.846016
Rwpos107_22 in107 sp22 11140.846016
Rwpos107_23 in107 sp23 3183.098862
Rwpos107_24 in107 sp24 3183.098862
Rwpos107_25 in107 sp25 3183.098862
Rwpos107_26 in107 sp26 11140.846016
Rwpos107_27 in107 sp27 11140.846016
Rwpos107_28 in107 sp28 3183.098862
Rwpos107_29 in107 sp29 3183.098862
Rwpos107_30 in107 sp30 3183.098862
Rwpos107_31 in107 sp31 3183.098862
Rwpos107_32 in107 sp32 11140.846016
Rwpos107_33 in107 sp33 11140.846016
Rwpos107_34 in107 sp34 11140.846016
Rwpos107_35 in107 sp35 3183.098862
Rwpos107_36 in107 sp36 3183.098862
Rwpos107_37 in107 sp37 3183.098862
Rwpos107_38 in107 sp38 3183.098862
Rwpos107_39 in107 sp39 3183.098862
Rwpos107_40 in107 sp40 3183.098862
Rwpos107_41 in107 sp41 3183.098862
Rwpos107_42 in107 sp42 11140.846016
Rwpos107_43 in107 sp43 11140.846016
Rwpos107_44 in107 sp44 11140.846016
Rwpos107_45 in107 sp45 3183.098862
Rwpos107_46 in107 sp46 3183.098862
Rwpos107_47 in107 sp47 3183.098862
Rwpos107_48 in107 sp48 11140.846016
Rwpos107_49 in107 sp49 11140.846016
Rwpos107_50 in107 sp50 11140.846016
Rwpos107_51 in107 sp51 11140.846016
Rwpos107_52 in107 sp52 11140.846016
Rwpos107_53 in107 sp53 11140.846016
Rwpos107_54 in107 sp54 11140.846016
Rwpos107_55 in107 sp55 3183.098862
Rwpos107_56 in107 sp56 11140.846016
Rwpos107_57 in107 sp57 3183.098862
Rwpos107_58 in107 sp58 11140.846016
Rwpos107_59 in107 sp59 11140.846016
Rwpos107_60 in107 sp60 3183.098862
Rwpos107_61 in107 sp61 3183.098862
Rwpos107_62 in107 sp62 3183.098862
Rwpos107_63 in107 sp63 11140.846016
Rwpos107_64 in107 sp64 11140.846016
Rwpos107_65 in107 sp65 11140.846016
Rwpos107_66 in107 sp66 11140.846016
Rwpos107_67 in107 sp67 3183.098862
Rwpos107_68 in107 sp68 11140.846016
Rwpos107_69 in107 sp69 3183.098862
Rwpos107_70 in107 sp70 11140.846016
Rwpos107_71 in107 sp71 3183.098862
Rwpos107_72 in107 sp72 11140.846016
Rwpos107_73 in107 sp73 11140.846016
Rwpos107_74 in107 sp74 3183.098862
Rwpos107_75 in107 sp75 11140.846016
Rwpos107_76 in107 sp76 3183.098862
Rwpos107_77 in107 sp77 11140.846016
Rwpos107_78 in107 sp78 3183.098862
Rwpos107_79 in107 sp79 3183.098862
Rwpos107_80 in107 sp80 3183.098862
Rwpos107_81 in107 sp81 11140.846016
Rwpos107_82 in107 sp82 11140.846016
Rwpos107_83 in107 sp83 11140.846016
Rwpos107_84 in107 sp84 11140.846016
Rwpos107_85 in107 sp85 11140.846016
Rwpos107_86 in107 sp86 11140.846016
Rwpos107_87 in107 sp87 3183.098862
Rwpos107_88 in107 sp88 3183.098862
Rwpos107_89 in107 sp89 3183.098862
Rwpos107_90 in107 sp90 11140.846016
Rwpos107_91 in107 sp91 11140.846016
Rwpos107_92 in107 sp92 11140.846016
Rwpos107_93 in107 sp93 11140.846016
Rwpos107_94 in107 sp94 11140.846016
Rwpos107_95 in107 sp95 3183.098862
Rwpos107_96 in107 sp96 11140.846016
Rwpos107_97 in107 sp97 11140.846016
Rwpos107_98 in107 sp98 11140.846016
Rwpos107_99 in107 sp99 3183.098862
Rwpos107_100 in107 sp100 11140.846016
Rwpos108_1 in108 sp1 3183.098862
Rwpos108_2 in108 sp2 3183.098862
Rwpos108_3 in108 sp3 11140.846016
Rwpos108_4 in108 sp4 11140.846016
Rwpos108_5 in108 sp5 3183.098862
Rwpos108_6 in108 sp6 3183.098862
Rwpos108_7 in108 sp7 3183.098862
Rwpos108_8 in108 sp8 3183.098862
Rwpos108_9 in108 sp9 3183.098862
Rwpos108_10 in108 sp10 3183.098862
Rwpos108_11 in108 sp11 11140.846016
Rwpos108_12 in108 sp12 3183.098862
Rwpos108_13 in108 sp13 11140.846016
Rwpos108_14 in108 sp14 11140.846016
Rwpos108_15 in108 sp15 3183.098862
Rwpos108_16 in108 sp16 3183.098862
Rwpos108_17 in108 sp17 11140.846016
Rwpos108_18 in108 sp18 11140.846016
Rwpos108_19 in108 sp19 11140.846016
Rwpos108_20 in108 sp20 11140.846016
Rwpos108_21 in108 sp21 3183.098862
Rwpos108_22 in108 sp22 3183.098862
Rwpos108_23 in108 sp23 3183.098862
Rwpos108_24 in108 sp24 11140.846016
Rwpos108_25 in108 sp25 3183.098862
Rwpos108_26 in108 sp26 3183.098862
Rwpos108_27 in108 sp27 3183.098862
Rwpos108_28 in108 sp28 11140.846016
Rwpos108_29 in108 sp29 3183.098862
Rwpos108_30 in108 sp30 3183.098862
Rwpos108_31 in108 sp31 3183.098862
Rwpos108_32 in108 sp32 11140.846016
Rwpos108_33 in108 sp33 3183.098862
Rwpos108_34 in108 sp34 11140.846016
Rwpos108_35 in108 sp35 3183.098862
Rwpos108_36 in108 sp36 3183.098862
Rwpos108_37 in108 sp37 3183.098862
Rwpos108_38 in108 sp38 3183.098862
Rwpos108_39 in108 sp39 3183.098862
Rwpos108_40 in108 sp40 11140.846016
Rwpos108_41 in108 sp41 11140.846016
Rwpos108_42 in108 sp42 3183.098862
Rwpos108_43 in108 sp43 11140.846016
Rwpos108_44 in108 sp44 3183.098862
Rwpos108_45 in108 sp45 3183.098862
Rwpos108_46 in108 sp46 11140.846016
Rwpos108_47 in108 sp47 11140.846016
Rwpos108_48 in108 sp48 3183.098862
Rwpos108_49 in108 sp49 3183.098862
Rwpos108_50 in108 sp50 3183.098862
Rwpos108_51 in108 sp51 3183.098862
Rwpos108_52 in108 sp52 11140.846016
Rwpos108_53 in108 sp53 3183.098862
Rwpos108_54 in108 sp54 11140.846016
Rwpos108_55 in108 sp55 11140.846016
Rwpos108_56 in108 sp56 3183.098862
Rwpos108_57 in108 sp57 3183.098862
Rwpos108_58 in108 sp58 3183.098862
Rwpos108_59 in108 sp59 11140.846016
Rwpos108_60 in108 sp60 11140.846016
Rwpos108_61 in108 sp61 3183.098862
Rwpos108_62 in108 sp62 11140.846016
Rwpos108_63 in108 sp63 11140.846016
Rwpos108_64 in108 sp64 3183.098862
Rwpos108_65 in108 sp65 11140.846016
Rwpos108_66 in108 sp66 11140.846016
Rwpos108_67 in108 sp67 3183.098862
Rwpos108_68 in108 sp68 11140.846016
Rwpos108_69 in108 sp69 3183.098862
Rwpos108_70 in108 sp70 11140.846016
Rwpos108_71 in108 sp71 3183.098862
Rwpos108_72 in108 sp72 3183.098862
Rwpos108_73 in108 sp73 3183.098862
Rwpos108_74 in108 sp74 11140.846016
Rwpos108_75 in108 sp75 11140.846016
Rwpos108_76 in108 sp76 3183.098862
Rwpos108_77 in108 sp77 3183.098862
Rwpos108_78 in108 sp78 11140.846016
Rwpos108_79 in108 sp79 3183.098862
Rwpos108_80 in108 sp80 11140.846016
Rwpos108_81 in108 sp81 3183.098862
Rwpos108_82 in108 sp82 11140.846016
Rwpos108_83 in108 sp83 11140.846016
Rwpos108_84 in108 sp84 11140.846016
Rwpos108_85 in108 sp85 3183.098862
Rwpos108_86 in108 sp86 3183.098862
Rwpos108_87 in108 sp87 11140.846016
Rwpos108_88 in108 sp88 3183.098862
Rwpos108_89 in108 sp89 11140.846016
Rwpos108_90 in108 sp90 11140.846016
Rwpos108_91 in108 sp91 3183.098862
Rwpos108_92 in108 sp92 11140.846016
Rwpos108_93 in108 sp93 11140.846016
Rwpos108_94 in108 sp94 3183.098862
Rwpos108_95 in108 sp95 11140.846016
Rwpos108_96 in108 sp96 11140.846016
Rwpos108_97 in108 sp97 3183.098862
Rwpos108_98 in108 sp98 11140.846016
Rwpos108_99 in108 sp99 3183.098862
Rwpos108_100 in108 sp100 11140.846016
Rwpos109_1 in109 sp1 11140.846016
Rwpos109_2 in109 sp2 11140.846016
Rwpos109_3 in109 sp3 11140.846016
Rwpos109_4 in109 sp4 11140.846016
Rwpos109_5 in109 sp5 3183.098862
Rwpos109_6 in109 sp6 3183.098862
Rwpos109_7 in109 sp7 3183.098862
Rwpos109_8 in109 sp8 3183.098862
Rwpos109_9 in109 sp9 11140.846016
Rwpos109_10 in109 sp10 3183.098862
Rwpos109_11 in109 sp11 3183.098862
Rwpos109_12 in109 sp12 3183.098862
Rwpos109_13 in109 sp13 11140.846016
Rwpos109_14 in109 sp14 11140.846016
Rwpos109_15 in109 sp15 3183.098862
Rwpos109_16 in109 sp16 3183.098862
Rwpos109_17 in109 sp17 11140.846016
Rwpos109_18 in109 sp18 11140.846016
Rwpos109_19 in109 sp19 11140.846016
Rwpos109_20 in109 sp20 11140.846016
Rwpos109_21 in109 sp21 3183.098862
Rwpos109_22 in109 sp22 11140.846016
Rwpos109_23 in109 sp23 11140.846016
Rwpos109_24 in109 sp24 11140.846016
Rwpos109_25 in109 sp25 3183.098862
Rwpos109_26 in109 sp26 3183.098862
Rwpos109_27 in109 sp27 3183.098862
Rwpos109_28 in109 sp28 11140.846016
Rwpos109_29 in109 sp29 11140.846016
Rwpos109_30 in109 sp30 11140.846016
Rwpos109_31 in109 sp31 3183.098862
Rwpos109_32 in109 sp32 3183.098862
Rwpos109_33 in109 sp33 11140.846016
Rwpos109_34 in109 sp34 3183.098862
Rwpos109_35 in109 sp35 3183.098862
Rwpos109_36 in109 sp36 11140.846016
Rwpos109_37 in109 sp37 11140.846016
Rwpos109_38 in109 sp38 3183.098862
Rwpos109_39 in109 sp39 3183.098862
Rwpos109_40 in109 sp40 3183.098862
Rwpos109_41 in109 sp41 11140.846016
Rwpos109_42 in109 sp42 11140.846016
Rwpos109_43 in109 sp43 11140.846016
Rwpos109_44 in109 sp44 3183.098862
Rwpos109_45 in109 sp45 3183.098862
Rwpos109_46 in109 sp46 3183.098862
Rwpos109_47 in109 sp47 11140.846016
Rwpos109_48 in109 sp48 11140.846016
Rwpos109_49 in109 sp49 11140.846016
Rwpos109_50 in109 sp50 11140.846016
Rwpos109_51 in109 sp51 11140.846016
Rwpos109_52 in109 sp52 11140.846016
Rwpos109_53 in109 sp53 3183.098862
Rwpos109_54 in109 sp54 11140.846016
Rwpos109_55 in109 sp55 11140.846016
Rwpos109_56 in109 sp56 3183.098862
Rwpos109_57 in109 sp57 3183.098862
Rwpos109_58 in109 sp58 11140.846016
Rwpos109_59 in109 sp59 11140.846016
Rwpos109_60 in109 sp60 3183.098862
Rwpos109_61 in109 sp61 3183.098862
Rwpos109_62 in109 sp62 3183.098862
Rwpos109_63 in109 sp63 11140.846016
Rwpos109_64 in109 sp64 11140.846016
Rwpos109_65 in109 sp65 11140.846016
Rwpos109_66 in109 sp66 3183.098862
Rwpos109_67 in109 sp67 11140.846016
Rwpos109_68 in109 sp68 3183.098862
Rwpos109_69 in109 sp69 11140.846016
Rwpos109_70 in109 sp70 11140.846016
Rwpos109_71 in109 sp71 3183.098862
Rwpos109_72 in109 sp72 3183.098862
Rwpos109_73 in109 sp73 11140.846016
Rwpos109_74 in109 sp74 11140.846016
Rwpos109_75 in109 sp75 11140.846016
Rwpos109_76 in109 sp76 3183.098862
Rwpos109_77 in109 sp77 3183.098862
Rwpos109_78 in109 sp78 3183.098862
Rwpos109_79 in109 sp79 3183.098862
Rwpos109_80 in109 sp80 3183.098862
Rwpos109_81 in109 sp81 11140.846016
Rwpos109_82 in109 sp82 3183.098862
Rwpos109_83 in109 sp83 3183.098862
Rwpos109_84 in109 sp84 11140.846016
Rwpos109_85 in109 sp85 3183.098862
Rwpos109_86 in109 sp86 11140.846016
Rwpos109_87 in109 sp87 3183.098862
Rwpos109_88 in109 sp88 11140.846016
Rwpos109_89 in109 sp89 3183.098862
Rwpos109_90 in109 sp90 11140.846016
Rwpos109_91 in109 sp91 11140.846016
Rwpos109_92 in109 sp92 3183.098862
Rwpos109_93 in109 sp93 3183.098862
Rwpos109_94 in109 sp94 3183.098862
Rwpos109_95 in109 sp95 11140.846016
Rwpos109_96 in109 sp96 11140.846016
Rwpos109_97 in109 sp97 11140.846016
Rwpos109_98 in109 sp98 11140.846016
Rwpos109_99 in109 sp99 11140.846016
Rwpos109_100 in109 sp100 3183.098862
Rwpos110_1 in110 sp1 11140.846016
Rwpos110_2 in110 sp2 11140.846016
Rwpos110_3 in110 sp3 11140.846016
Rwpos110_4 in110 sp4 11140.846016
Rwpos110_5 in110 sp5 11140.846016
Rwpos110_6 in110 sp6 3183.098862
Rwpos110_7 in110 sp7 3183.098862
Rwpos110_8 in110 sp8 3183.098862
Rwpos110_9 in110 sp9 11140.846016
Rwpos110_10 in110 sp10 3183.098862
Rwpos110_11 in110 sp11 11140.846016
Rwpos110_12 in110 sp12 3183.098862
Rwpos110_13 in110 sp13 11140.846016
Rwpos110_14 in110 sp14 3183.098862
Rwpos110_15 in110 sp15 3183.098862
Rwpos110_16 in110 sp16 11140.846016
Rwpos110_17 in110 sp17 11140.846016
Rwpos110_18 in110 sp18 11140.846016
Rwpos110_19 in110 sp19 3183.098862
Rwpos110_20 in110 sp20 3183.098862
Rwpos110_21 in110 sp21 11140.846016
Rwpos110_22 in110 sp22 3183.098862
Rwpos110_23 in110 sp23 3183.098862
Rwpos110_24 in110 sp24 3183.098862
Rwpos110_25 in110 sp25 3183.098862
Rwpos110_26 in110 sp26 3183.098862
Rwpos110_27 in110 sp27 3183.098862
Rwpos110_28 in110 sp28 3183.098862
Rwpos110_29 in110 sp29 11140.846016
Rwpos110_30 in110 sp30 3183.098862
Rwpos110_31 in110 sp31 3183.098862
Rwpos110_32 in110 sp32 3183.098862
Rwpos110_33 in110 sp33 3183.098862
Rwpos110_34 in110 sp34 11140.846016
Rwpos110_35 in110 sp35 3183.098862
Rwpos110_36 in110 sp36 3183.098862
Rwpos110_37 in110 sp37 3183.098862
Rwpos110_38 in110 sp38 3183.098862
Rwpos110_39 in110 sp39 3183.098862
Rwpos110_40 in110 sp40 11140.846016
Rwpos110_41 in110 sp41 11140.846016
Rwpos110_42 in110 sp42 3183.098862
Rwpos110_43 in110 sp43 3183.098862
Rwpos110_44 in110 sp44 3183.098862
Rwpos110_45 in110 sp45 3183.098862
Rwpos110_46 in110 sp46 3183.098862
Rwpos110_47 in110 sp47 3183.098862
Rwpos110_48 in110 sp48 3183.098862
Rwpos110_49 in110 sp49 11140.846016
Rwpos110_50 in110 sp50 11140.846016
Rwpos110_51 in110 sp51 11140.846016
Rwpos110_52 in110 sp52 3183.098862
Rwpos110_53 in110 sp53 3183.098862
Rwpos110_54 in110 sp54 3183.098862
Rwpos110_55 in110 sp55 3183.098862
Rwpos110_56 in110 sp56 3183.098862
Rwpos110_57 in110 sp57 3183.098862
Rwpos110_58 in110 sp58 11140.846016
Rwpos110_59 in110 sp59 11140.846016
Rwpos110_60 in110 sp60 3183.098862
Rwpos110_61 in110 sp61 11140.846016
Rwpos110_62 in110 sp62 3183.098862
Rwpos110_63 in110 sp63 11140.846016
Rwpos110_64 in110 sp64 3183.098862
Rwpos110_65 in110 sp65 3183.098862
Rwpos110_66 in110 sp66 11140.846016
Rwpos110_67 in110 sp67 3183.098862
Rwpos110_68 in110 sp68 3183.098862
Rwpos110_69 in110 sp69 3183.098862
Rwpos110_70 in110 sp70 3183.098862
Rwpos110_71 in110 sp71 11140.846016
Rwpos110_72 in110 sp72 11140.846016
Rwpos110_73 in110 sp73 11140.846016
Rwpos110_74 in110 sp74 3183.098862
Rwpos110_75 in110 sp75 3183.098862
Rwpos110_76 in110 sp76 3183.098862
Rwpos110_77 in110 sp77 11140.846016
Rwpos110_78 in110 sp78 3183.098862
Rwpos110_79 in110 sp79 3183.098862
Rwpos110_80 in110 sp80 11140.846016
Rwpos110_81 in110 sp81 11140.846016
Rwpos110_82 in110 sp82 3183.098862
Rwpos110_83 in110 sp83 3183.098862
Rwpos110_84 in110 sp84 3183.098862
Rwpos110_85 in110 sp85 11140.846016
Rwpos110_86 in110 sp86 3183.098862
Rwpos110_87 in110 sp87 3183.098862
Rwpos110_88 in110 sp88 3183.098862
Rwpos110_89 in110 sp89 11140.846016
Rwpos110_90 in110 sp90 11140.846016
Rwpos110_91 in110 sp91 3183.098862
Rwpos110_92 in110 sp92 3183.098862
Rwpos110_93 in110 sp93 11140.846016
Rwpos110_94 in110 sp94 3183.098862
Rwpos110_95 in110 sp95 11140.846016
Rwpos110_96 in110 sp96 3183.098862
Rwpos110_97 in110 sp97 11140.846016
Rwpos110_98 in110 sp98 3183.098862
Rwpos110_99 in110 sp99 3183.098862
Rwpos110_100 in110 sp100 11140.846016
Rwpos111_1 in111 sp1 3183.098862
Rwpos111_2 in111 sp2 3183.098862
Rwpos111_3 in111 sp3 3183.098862
Rwpos111_4 in111 sp4 3183.098862
Rwpos111_5 in111 sp5 11140.846016
Rwpos111_6 in111 sp6 3183.098862
Rwpos111_7 in111 sp7 3183.098862
Rwpos111_8 in111 sp8 3183.098862
Rwpos111_9 in111 sp9 11140.846016
Rwpos111_10 in111 sp10 3183.098862
Rwpos111_11 in111 sp11 11140.846016
Rwpos111_12 in111 sp12 3183.098862
Rwpos111_13 in111 sp13 3183.098862
Rwpos111_14 in111 sp14 3183.098862
Rwpos111_15 in111 sp15 3183.098862
Rwpos111_16 in111 sp16 3183.098862
Rwpos111_17 in111 sp17 3183.098862
Rwpos111_18 in111 sp18 3183.098862
Rwpos111_19 in111 sp19 3183.098862
Rwpos111_20 in111 sp20 3183.098862
Rwpos111_21 in111 sp21 11140.846016
Rwpos111_22 in111 sp22 11140.846016
Rwpos111_23 in111 sp23 11140.846016
Rwpos111_24 in111 sp24 3183.098862
Rwpos111_25 in111 sp25 3183.098862
Rwpos111_26 in111 sp26 3183.098862
Rwpos111_27 in111 sp27 11140.846016
Rwpos111_28 in111 sp28 11140.846016
Rwpos111_29 in111 sp29 11140.846016
Rwpos111_30 in111 sp30 3183.098862
Rwpos111_31 in111 sp31 3183.098862
Rwpos111_32 in111 sp32 3183.098862
Rwpos111_33 in111 sp33 3183.098862
Rwpos111_34 in111 sp34 3183.098862
Rwpos111_35 in111 sp35 11140.846016
Rwpos111_36 in111 sp36 11140.846016
Rwpos111_37 in111 sp37 11140.846016
Rwpos111_38 in111 sp38 11140.846016
Rwpos111_39 in111 sp39 3183.098862
Rwpos111_40 in111 sp40 3183.098862
Rwpos111_41 in111 sp41 3183.098862
Rwpos111_42 in111 sp42 3183.098862
Rwpos111_43 in111 sp43 11140.846016
Rwpos111_44 in111 sp44 3183.098862
Rwpos111_45 in111 sp45 11140.846016
Rwpos111_46 in111 sp46 3183.098862
Rwpos111_47 in111 sp47 11140.846016
Rwpos111_48 in111 sp48 11140.846016
Rwpos111_49 in111 sp49 3183.098862
Rwpos111_50 in111 sp50 3183.098862
Rwpos111_51 in111 sp51 3183.098862
Rwpos111_52 in111 sp52 3183.098862
Rwpos111_53 in111 sp53 3183.098862
Rwpos111_54 in111 sp54 11140.846016
Rwpos111_55 in111 sp55 11140.846016
Rwpos111_56 in111 sp56 3183.098862
Rwpos111_57 in111 sp57 3183.098862
Rwpos111_58 in111 sp58 3183.098862
Rwpos111_59 in111 sp59 11140.846016
Rwpos111_60 in111 sp60 3183.098862
Rwpos111_61 in111 sp61 11140.846016
Rwpos111_62 in111 sp62 3183.098862
Rwpos111_63 in111 sp63 11140.846016
Rwpos111_64 in111 sp64 11140.846016
Rwpos111_65 in111 sp65 3183.098862
Rwpos111_66 in111 sp66 3183.098862
Rwpos111_67 in111 sp67 3183.098862
Rwpos111_68 in111 sp68 3183.098862
Rwpos111_69 in111 sp69 3183.098862
Rwpos111_70 in111 sp70 3183.098862
Rwpos111_71 in111 sp71 11140.846016
Rwpos111_72 in111 sp72 3183.098862
Rwpos111_73 in111 sp73 11140.846016
Rwpos111_74 in111 sp74 3183.098862
Rwpos111_75 in111 sp75 11140.846016
Rwpos111_76 in111 sp76 3183.098862
Rwpos111_77 in111 sp77 11140.846016
Rwpos111_78 in111 sp78 3183.098862
Rwpos111_79 in111 sp79 11140.846016
Rwpos111_80 in111 sp80 11140.846016
Rwpos111_81 in111 sp81 11140.846016
Rwpos111_82 in111 sp82 11140.846016
Rwpos111_83 in111 sp83 3183.098862
Rwpos111_84 in111 sp84 11140.846016
Rwpos111_85 in111 sp85 11140.846016
Rwpos111_86 in111 sp86 11140.846016
Rwpos111_87 in111 sp87 11140.846016
Rwpos111_88 in111 sp88 3183.098862
Rwpos111_89 in111 sp89 3183.098862
Rwpos111_90 in111 sp90 11140.846016
Rwpos111_91 in111 sp91 11140.846016
Rwpos111_92 in111 sp92 3183.098862
Rwpos111_93 in111 sp93 11140.846016
Rwpos111_94 in111 sp94 3183.098862
Rwpos111_95 in111 sp95 11140.846016
Rwpos111_96 in111 sp96 11140.846016
Rwpos111_97 in111 sp97 11140.846016
Rwpos111_98 in111 sp98 3183.098862
Rwpos111_99 in111 sp99 3183.098862
Rwpos111_100 in111 sp100 3183.098862
Rwpos112_1 in112 sp1 3183.098862
Rwpos112_2 in112 sp2 3183.098862
Rwpos112_3 in112 sp3 11140.846016
Rwpos112_4 in112 sp4 11140.846016
Rwpos112_5 in112 sp5 11140.846016
Rwpos112_6 in112 sp6 3183.098862
Rwpos112_7 in112 sp7 11140.846016
Rwpos112_8 in112 sp8 11140.846016
Rwpos112_9 in112 sp9 3183.098862
Rwpos112_10 in112 sp10 3183.098862
Rwpos112_11 in112 sp11 11140.846016
Rwpos112_12 in112 sp12 3183.098862
Rwpos112_13 in112 sp13 11140.846016
Rwpos112_14 in112 sp14 3183.098862
Rwpos112_15 in112 sp15 3183.098862
Rwpos112_16 in112 sp16 11140.846016
Rwpos112_17 in112 sp17 11140.846016
Rwpos112_18 in112 sp18 11140.846016
Rwpos112_19 in112 sp19 3183.098862
Rwpos112_20 in112 sp20 3183.098862
Rwpos112_21 in112 sp21 11140.846016
Rwpos112_22 in112 sp22 3183.098862
Rwpos112_23 in112 sp23 11140.846016
Rwpos112_24 in112 sp24 3183.098862
Rwpos112_25 in112 sp25 3183.098862
Rwpos112_26 in112 sp26 3183.098862
Rwpos112_27 in112 sp27 3183.098862
Rwpos112_28 in112 sp28 11140.846016
Rwpos112_29 in112 sp29 11140.846016
Rwpos112_30 in112 sp30 3183.098862
Rwpos112_31 in112 sp31 3183.098862
Rwpos112_32 in112 sp32 3183.098862
Rwpos112_33 in112 sp33 11140.846016
Rwpos112_34 in112 sp34 3183.098862
Rwpos112_35 in112 sp35 3183.098862
Rwpos112_36 in112 sp36 11140.846016
Rwpos112_37 in112 sp37 11140.846016
Rwpos112_38 in112 sp38 11140.846016
Rwpos112_39 in112 sp39 11140.846016
Rwpos112_40 in112 sp40 11140.846016
Rwpos112_41 in112 sp41 3183.098862
Rwpos112_42 in112 sp42 11140.846016
Rwpos112_43 in112 sp43 3183.098862
Rwpos112_44 in112 sp44 3183.098862
Rwpos112_45 in112 sp45 11140.846016
Rwpos112_46 in112 sp46 11140.846016
Rwpos112_47 in112 sp47 11140.846016
Rwpos112_48 in112 sp48 11140.846016
Rwpos112_49 in112 sp49 3183.098862
Rwpos112_50 in112 sp50 11140.846016
Rwpos112_51 in112 sp51 3183.098862
Rwpos112_52 in112 sp52 11140.846016
Rwpos112_53 in112 sp53 11140.846016
Rwpos112_54 in112 sp54 11140.846016
Rwpos112_55 in112 sp55 11140.846016
Rwpos112_56 in112 sp56 3183.098862
Rwpos112_57 in112 sp57 3183.098862
Rwpos112_58 in112 sp58 3183.098862
Rwpos112_59 in112 sp59 11140.846016
Rwpos112_60 in112 sp60 11140.846016
Rwpos112_61 in112 sp61 11140.846016
Rwpos112_62 in112 sp62 3183.098862
Rwpos112_63 in112 sp63 3183.098862
Rwpos112_64 in112 sp64 3183.098862
Rwpos112_65 in112 sp65 3183.098862
Rwpos112_66 in112 sp66 11140.846016
Rwpos112_67 in112 sp67 3183.098862
Rwpos112_68 in112 sp68 11140.846016
Rwpos112_69 in112 sp69 11140.846016
Rwpos112_70 in112 sp70 11140.846016
Rwpos112_71 in112 sp71 11140.846016
Rwpos112_72 in112 sp72 3183.098862
Rwpos112_73 in112 sp73 11140.846016
Rwpos112_74 in112 sp74 11140.846016
Rwpos112_75 in112 sp75 11140.846016
Rwpos112_76 in112 sp76 11140.846016
Rwpos112_77 in112 sp77 11140.846016
Rwpos112_78 in112 sp78 11140.846016
Rwpos112_79 in112 sp79 11140.846016
Rwpos112_80 in112 sp80 3183.098862
Rwpos112_81 in112 sp81 3183.098862
Rwpos112_82 in112 sp82 3183.098862
Rwpos112_83 in112 sp83 3183.098862
Rwpos112_84 in112 sp84 3183.098862
Rwpos112_85 in112 sp85 3183.098862
Rwpos112_86 in112 sp86 3183.098862
Rwpos112_87 in112 sp87 11140.846016
Rwpos112_88 in112 sp88 11140.846016
Rwpos112_89 in112 sp89 3183.098862
Rwpos112_90 in112 sp90 11140.846016
Rwpos112_91 in112 sp91 3183.098862
Rwpos112_92 in112 sp92 3183.098862
Rwpos112_93 in112 sp93 3183.098862
Rwpos112_94 in112 sp94 11140.846016
Rwpos112_95 in112 sp95 11140.846016
Rwpos112_96 in112 sp96 11140.846016
Rwpos112_97 in112 sp97 3183.098862
Rwpos112_98 in112 sp98 3183.098862
Rwpos112_99 in112 sp99 3183.098862
Rwpos112_100 in112 sp100 3183.098862
Rwpos113_1 in113 sp1 3183.098862
Rwpos113_2 in113 sp2 3183.098862
Rwpos113_3 in113 sp3 11140.846016
Rwpos113_4 in113 sp4 11140.846016
Rwpos113_5 in113 sp5 11140.846016
Rwpos113_6 in113 sp6 11140.846016
Rwpos113_7 in113 sp7 3183.098862
Rwpos113_8 in113 sp8 3183.098862
Rwpos113_9 in113 sp9 3183.098862
Rwpos113_10 in113 sp10 3183.098862
Rwpos113_11 in113 sp11 3183.098862
Rwpos113_12 in113 sp12 11140.846016
Rwpos113_13 in113 sp13 3183.098862
Rwpos113_14 in113 sp14 11140.846016
Rwpos113_15 in113 sp15 11140.846016
Rwpos113_16 in113 sp16 11140.846016
Rwpos113_17 in113 sp17 11140.846016
Rwpos113_18 in113 sp18 3183.098862
Rwpos113_19 in113 sp19 11140.846016
Rwpos113_20 in113 sp20 3183.098862
Rwpos113_21 in113 sp21 3183.098862
Rwpos113_22 in113 sp22 11140.846016
Rwpos113_23 in113 sp23 11140.846016
Rwpos113_24 in113 sp24 3183.098862
Rwpos113_25 in113 sp25 11140.846016
Rwpos113_26 in113 sp26 11140.846016
Rwpos113_27 in113 sp27 3183.098862
Rwpos113_28 in113 sp28 11140.846016
Rwpos113_29 in113 sp29 3183.098862
Rwpos113_30 in113 sp30 11140.846016
Rwpos113_31 in113 sp31 11140.846016
Rwpos113_32 in113 sp32 11140.846016
Rwpos113_33 in113 sp33 11140.846016
Rwpos113_34 in113 sp34 3183.098862
Rwpos113_35 in113 sp35 3183.098862
Rwpos113_36 in113 sp36 11140.846016
Rwpos113_37 in113 sp37 11140.846016
Rwpos113_38 in113 sp38 11140.846016
Rwpos113_39 in113 sp39 11140.846016
Rwpos113_40 in113 sp40 11140.846016
Rwpos113_41 in113 sp41 3183.098862
Rwpos113_42 in113 sp42 3183.098862
Rwpos113_43 in113 sp43 3183.098862
Rwpos113_44 in113 sp44 11140.846016
Rwpos113_45 in113 sp45 11140.846016
Rwpos113_46 in113 sp46 11140.846016
Rwpos113_47 in113 sp47 11140.846016
Rwpos113_48 in113 sp48 11140.846016
Rwpos113_49 in113 sp49 11140.846016
Rwpos113_50 in113 sp50 11140.846016
Rwpos113_51 in113 sp51 11140.846016
Rwpos113_52 in113 sp52 3183.098862
Rwpos113_53 in113 sp53 3183.098862
Rwpos113_54 in113 sp54 3183.098862
Rwpos113_55 in113 sp55 11140.846016
Rwpos113_56 in113 sp56 11140.846016
Rwpos113_57 in113 sp57 11140.846016
Rwpos113_58 in113 sp58 11140.846016
Rwpos113_59 in113 sp59 3183.098862
Rwpos113_60 in113 sp60 3183.098862
Rwpos113_61 in113 sp61 11140.846016
Rwpos113_62 in113 sp62 3183.098862
Rwpos113_63 in113 sp63 11140.846016
Rwpos113_64 in113 sp64 3183.098862
Rwpos113_65 in113 sp65 3183.098862
Rwpos113_66 in113 sp66 11140.846016
Rwpos113_67 in113 sp67 11140.846016
Rwpos113_68 in113 sp68 11140.846016
Rwpos113_69 in113 sp69 11140.846016
Rwpos113_70 in113 sp70 3183.098862
Rwpos113_71 in113 sp71 3183.098862
Rwpos113_72 in113 sp72 11140.846016
Rwpos113_73 in113 sp73 11140.846016
Rwpos113_74 in113 sp74 3183.098862
Rwpos113_75 in113 sp75 11140.846016
Rwpos113_76 in113 sp76 3183.098862
Rwpos113_77 in113 sp77 11140.846016
Rwpos113_78 in113 sp78 3183.098862
Rwpos113_79 in113 sp79 11140.846016
Rwpos113_80 in113 sp80 11140.846016
Rwpos113_81 in113 sp81 11140.846016
Rwpos113_82 in113 sp82 11140.846016
Rwpos113_83 in113 sp83 11140.846016
Rwpos113_84 in113 sp84 11140.846016
Rwpos113_85 in113 sp85 11140.846016
Rwpos113_86 in113 sp86 3183.098862
Rwpos113_87 in113 sp87 3183.098862
Rwpos113_88 in113 sp88 3183.098862
Rwpos113_89 in113 sp89 11140.846016
Rwpos113_90 in113 sp90 3183.098862
Rwpos113_91 in113 sp91 3183.098862
Rwpos113_92 in113 sp92 3183.098862
Rwpos113_93 in113 sp93 3183.098862
Rwpos113_94 in113 sp94 11140.846016
Rwpos113_95 in113 sp95 11140.846016
Rwpos113_96 in113 sp96 11140.846016
Rwpos113_97 in113 sp97 11140.846016
Rwpos113_98 in113 sp98 3183.098862
Rwpos113_99 in113 sp99 11140.846016
Rwpos113_100 in113 sp100 3183.098862
Rwpos114_1 in114 sp1 3183.098862
Rwpos114_2 in114 sp2 3183.098862
Rwpos114_3 in114 sp3 11140.846016
Rwpos114_4 in114 sp4 3183.098862
Rwpos114_5 in114 sp5 11140.846016
Rwpos114_6 in114 sp6 3183.098862
Rwpos114_7 in114 sp7 3183.098862
Rwpos114_8 in114 sp8 3183.098862
Rwpos114_9 in114 sp9 3183.098862
Rwpos114_10 in114 sp10 11140.846016
Rwpos114_11 in114 sp11 11140.846016
Rwpos114_12 in114 sp12 3183.098862
Rwpos114_13 in114 sp13 11140.846016
Rwpos114_14 in114 sp14 3183.098862
Rwpos114_15 in114 sp15 11140.846016
Rwpos114_16 in114 sp16 3183.098862
Rwpos114_17 in114 sp17 3183.098862
Rwpos114_18 in114 sp18 11140.846016
Rwpos114_19 in114 sp19 3183.098862
Rwpos114_20 in114 sp20 3183.098862
Rwpos114_21 in114 sp21 11140.846016
Rwpos114_22 in114 sp22 3183.098862
Rwpos114_23 in114 sp23 11140.846016
Rwpos114_24 in114 sp24 11140.846016
Rwpos114_25 in114 sp25 3183.098862
Rwpos114_26 in114 sp26 3183.098862
Rwpos114_27 in114 sp27 3183.098862
Rwpos114_28 in114 sp28 3183.098862
Rwpos114_29 in114 sp29 11140.846016
Rwpos114_30 in114 sp30 3183.098862
Rwpos114_31 in114 sp31 11140.846016
Rwpos114_32 in114 sp32 11140.846016
Rwpos114_33 in114 sp33 11140.846016
Rwpos114_34 in114 sp34 11140.846016
Rwpos114_35 in114 sp35 3183.098862
Rwpos114_36 in114 sp36 11140.846016
Rwpos114_37 in114 sp37 3183.098862
Rwpos114_38 in114 sp38 3183.098862
Rwpos114_39 in114 sp39 3183.098862
Rwpos114_40 in114 sp40 3183.098862
Rwpos114_41 in114 sp41 3183.098862
Rwpos114_42 in114 sp42 3183.098862
Rwpos114_43 in114 sp43 11140.846016
Rwpos114_44 in114 sp44 3183.098862
Rwpos114_45 in114 sp45 11140.846016
Rwpos114_46 in114 sp46 3183.098862
Rwpos114_47 in114 sp47 11140.846016
Rwpos114_48 in114 sp48 11140.846016
Rwpos114_49 in114 sp49 11140.846016
Rwpos114_50 in114 sp50 3183.098862
Rwpos114_51 in114 sp51 3183.098862
Rwpos114_52 in114 sp52 11140.846016
Rwpos114_53 in114 sp53 3183.098862
Rwpos114_54 in114 sp54 3183.098862
Rwpos114_55 in114 sp55 11140.846016
Rwpos114_56 in114 sp56 3183.098862
Rwpos114_57 in114 sp57 3183.098862
Rwpos114_58 in114 sp58 3183.098862
Rwpos114_59 in114 sp59 11140.846016
Rwpos114_60 in114 sp60 3183.098862
Rwpos114_61 in114 sp61 11140.846016
Rwpos114_62 in114 sp62 3183.098862
Rwpos114_63 in114 sp63 11140.846016
Rwpos114_64 in114 sp64 11140.846016
Rwpos114_65 in114 sp65 11140.846016
Rwpos114_66 in114 sp66 11140.846016
Rwpos114_67 in114 sp67 3183.098862
Rwpos114_68 in114 sp68 11140.846016
Rwpos114_69 in114 sp69 3183.098862
Rwpos114_70 in114 sp70 3183.098862
Rwpos114_71 in114 sp71 3183.098862
Rwpos114_72 in114 sp72 3183.098862
Rwpos114_73 in114 sp73 3183.098862
Rwpos114_74 in114 sp74 3183.098862
Rwpos114_75 in114 sp75 11140.846016
Rwpos114_76 in114 sp76 3183.098862
Rwpos114_77 in114 sp77 11140.846016
Rwpos114_78 in114 sp78 3183.098862
Rwpos114_79 in114 sp79 11140.846016
Rwpos114_80 in114 sp80 11140.846016
Rwpos114_81 in114 sp81 11140.846016
Rwpos114_82 in114 sp82 3183.098862
Rwpos114_83 in114 sp83 3183.098862
Rwpos114_84 in114 sp84 3183.098862
Rwpos114_85 in114 sp85 11140.846016
Rwpos114_86 in114 sp86 3183.098862
Rwpos114_87 in114 sp87 11140.846016
Rwpos114_88 in114 sp88 3183.098862
Rwpos114_89 in114 sp89 3183.098862
Rwpos114_90 in114 sp90 3183.098862
Rwpos114_91 in114 sp91 11140.846016
Rwpos114_92 in114 sp92 3183.098862
Rwpos114_93 in114 sp93 11140.846016
Rwpos114_94 in114 sp94 3183.098862
Rwpos114_95 in114 sp95 11140.846016
Rwpos114_96 in114 sp96 11140.846016
Rwpos114_97 in114 sp97 11140.846016
Rwpos114_98 in114 sp98 3183.098862
Rwpos114_99 in114 sp99 3183.098862
Rwpos114_100 in114 sp100 11140.846016
Rwpos115_1 in115 sp1 3183.098862
Rwpos115_2 in115 sp2 3183.098862
Rwpos115_3 in115 sp3 11140.846016
Rwpos115_4 in115 sp4 3183.098862
Rwpos115_5 in115 sp5 3183.098862
Rwpos115_6 in115 sp6 3183.098862
Rwpos115_7 in115 sp7 11140.846016
Rwpos115_8 in115 sp8 11140.846016
Rwpos115_9 in115 sp9 11140.846016
Rwpos115_10 in115 sp10 3183.098862
Rwpos115_11 in115 sp11 11140.846016
Rwpos115_12 in115 sp12 11140.846016
Rwpos115_13 in115 sp13 11140.846016
Rwpos115_14 in115 sp14 3183.098862
Rwpos115_15 in115 sp15 3183.098862
Rwpos115_16 in115 sp16 11140.846016
Rwpos115_17 in115 sp17 3183.098862
Rwpos115_18 in115 sp18 3183.098862
Rwpos115_19 in115 sp19 11140.846016
Rwpos115_20 in115 sp20 3183.098862
Rwpos115_21 in115 sp21 3183.098862
Rwpos115_22 in115 sp22 3183.098862
Rwpos115_23 in115 sp23 11140.846016
Rwpos115_24 in115 sp24 3183.098862
Rwpos115_25 in115 sp25 11140.846016
Rwpos115_26 in115 sp26 3183.098862
Rwpos115_27 in115 sp27 11140.846016
Rwpos115_28 in115 sp28 3183.098862
Rwpos115_29 in115 sp29 3183.098862
Rwpos115_30 in115 sp30 3183.098862
Rwpos115_31 in115 sp31 3183.098862
Rwpos115_32 in115 sp32 3183.098862
Rwpos115_33 in115 sp33 3183.098862
Rwpos115_34 in115 sp34 3183.098862
Rwpos115_35 in115 sp35 3183.098862
Rwpos115_36 in115 sp36 3183.098862
Rwpos115_37 in115 sp37 3183.098862
Rwpos115_38 in115 sp38 3183.098862
Rwpos115_39 in115 sp39 11140.846016
Rwpos115_40 in115 sp40 3183.098862
Rwpos115_41 in115 sp41 11140.846016
Rwpos115_42 in115 sp42 3183.098862
Rwpos115_43 in115 sp43 11140.846016
Rwpos115_44 in115 sp44 3183.098862
Rwpos115_45 in115 sp45 11140.846016
Rwpos115_46 in115 sp46 3183.098862
Rwpos115_47 in115 sp47 3183.098862
Rwpos115_48 in115 sp48 3183.098862
Rwpos115_49 in115 sp49 3183.098862
Rwpos115_50 in115 sp50 3183.098862
Rwpos115_51 in115 sp51 3183.098862
Rwpos115_52 in115 sp52 11140.846016
Rwpos115_53 in115 sp53 3183.098862
Rwpos115_54 in115 sp54 3183.098862
Rwpos115_55 in115 sp55 11140.846016
Rwpos115_56 in115 sp56 3183.098862
Rwpos115_57 in115 sp57 11140.846016
Rwpos115_58 in115 sp58 3183.098862
Rwpos115_59 in115 sp59 11140.846016
Rwpos115_60 in115 sp60 11140.846016
Rwpos115_61 in115 sp61 11140.846016
Rwpos115_62 in115 sp62 3183.098862
Rwpos115_63 in115 sp63 3183.098862
Rwpos115_64 in115 sp64 3183.098862
Rwpos115_65 in115 sp65 11140.846016
Rwpos115_66 in115 sp66 3183.098862
Rwpos115_67 in115 sp67 3183.098862
Rwpos115_68 in115 sp68 3183.098862
Rwpos115_69 in115 sp69 3183.098862
Rwpos115_70 in115 sp70 3183.098862
Rwpos115_71 in115 sp71 11140.846016
Rwpos115_72 in115 sp72 3183.098862
Rwpos115_73 in115 sp73 3183.098862
Rwpos115_74 in115 sp74 3183.098862
Rwpos115_75 in115 sp75 11140.846016
Rwpos115_76 in115 sp76 3183.098862
Rwpos115_77 in115 sp77 11140.846016
Rwpos115_78 in115 sp78 3183.098862
Rwpos115_79 in115 sp79 11140.846016
Rwpos115_80 in115 sp80 11140.846016
Rwpos115_81 in115 sp81 11140.846016
Rwpos115_82 in115 sp82 3183.098862
Rwpos115_83 in115 sp83 3183.098862
Rwpos115_84 in115 sp84 3183.098862
Rwpos115_85 in115 sp85 3183.098862
Rwpos115_86 in115 sp86 3183.098862
Rwpos115_87 in115 sp87 11140.846016
Rwpos115_88 in115 sp88 3183.098862
Rwpos115_89 in115 sp89 11140.846016
Rwpos115_90 in115 sp90 3183.098862
Rwpos115_91 in115 sp91 11140.846016
Rwpos115_92 in115 sp92 3183.098862
Rwpos115_93 in115 sp93 3183.098862
Rwpos115_94 in115 sp94 3183.098862
Rwpos115_95 in115 sp95 3183.098862
Rwpos115_96 in115 sp96 3183.098862
Rwpos115_97 in115 sp97 3183.098862
Rwpos115_98 in115 sp98 3183.098862
Rwpos115_99 in115 sp99 11140.846016
Rwpos115_100 in115 sp100 3183.098862
Rwpos116_1 in116 sp1 11140.846016
Rwpos116_2 in116 sp2 11140.846016
Rwpos116_3 in116 sp3 3183.098862
Rwpos116_4 in116 sp4 11140.846016
Rwpos116_5 in116 sp5 11140.846016
Rwpos116_6 in116 sp6 3183.098862
Rwpos116_7 in116 sp7 11140.846016
Rwpos116_8 in116 sp8 11140.846016
Rwpos116_9 in116 sp9 3183.098862
Rwpos116_10 in116 sp10 3183.098862
Rwpos116_11 in116 sp11 3183.098862
Rwpos116_12 in116 sp12 3183.098862
Rwpos116_13 in116 sp13 3183.098862
Rwpos116_14 in116 sp14 3183.098862
Rwpos116_15 in116 sp15 3183.098862
Rwpos116_16 in116 sp16 3183.098862
Rwpos116_17 in116 sp17 3183.098862
Rwpos116_18 in116 sp18 3183.098862
Rwpos116_19 in116 sp19 3183.098862
Rwpos116_20 in116 sp20 3183.098862
Rwpos116_21 in116 sp21 3183.098862
Rwpos116_22 in116 sp22 3183.098862
Rwpos116_23 in116 sp23 11140.846016
Rwpos116_24 in116 sp24 3183.098862
Rwpos116_25 in116 sp25 11140.846016
Rwpos116_26 in116 sp26 11140.846016
Rwpos116_27 in116 sp27 3183.098862
Rwpos116_28 in116 sp28 11140.846016
Rwpos116_29 in116 sp29 11140.846016
Rwpos116_30 in116 sp30 3183.098862
Rwpos116_31 in116 sp31 11140.846016
Rwpos116_32 in116 sp32 11140.846016
Rwpos116_33 in116 sp33 3183.098862
Rwpos116_34 in116 sp34 11140.846016
Rwpos116_35 in116 sp35 3183.098862
Rwpos116_36 in116 sp36 11140.846016
Rwpos116_37 in116 sp37 3183.098862
Rwpos116_38 in116 sp38 3183.098862
Rwpos116_39 in116 sp39 11140.846016
Rwpos116_40 in116 sp40 11140.846016
Rwpos116_41 in116 sp41 3183.098862
Rwpos116_42 in116 sp42 3183.098862
Rwpos116_43 in116 sp43 3183.098862
Rwpos116_44 in116 sp44 3183.098862
Rwpos116_45 in116 sp45 3183.098862
Rwpos116_46 in116 sp46 3183.098862
Rwpos116_47 in116 sp47 11140.846016
Rwpos116_48 in116 sp48 3183.098862
Rwpos116_49 in116 sp49 11140.846016
Rwpos116_50 in116 sp50 3183.098862
Rwpos116_51 in116 sp51 11140.846016
Rwpos116_52 in116 sp52 11140.846016
Rwpos116_53 in116 sp53 3183.098862
Rwpos116_54 in116 sp54 3183.098862
Rwpos116_55 in116 sp55 3183.098862
Rwpos116_56 in116 sp56 11140.846016
Rwpos116_57 in116 sp57 3183.098862
Rwpos116_58 in116 sp58 11140.846016
Rwpos116_59 in116 sp59 3183.098862
Rwpos116_60 in116 sp60 11140.846016
Rwpos116_61 in116 sp61 11140.846016
Rwpos116_62 in116 sp62 11140.846016
Rwpos116_63 in116 sp63 3183.098862
Rwpos116_64 in116 sp64 3183.098862
Rwpos116_65 in116 sp65 3183.098862
Rwpos116_66 in116 sp66 3183.098862
Rwpos116_67 in116 sp67 11140.846016
Rwpos116_68 in116 sp68 11140.846016
Rwpos116_69 in116 sp69 11140.846016
Rwpos116_70 in116 sp70 11140.846016
Rwpos116_71 in116 sp71 3183.098862
Rwpos116_72 in116 sp72 3183.098862
Rwpos116_73 in116 sp73 3183.098862
Rwpos116_74 in116 sp74 3183.098862
Rwpos116_75 in116 sp75 3183.098862
Rwpos116_76 in116 sp76 3183.098862
Rwpos116_77 in116 sp77 3183.098862
Rwpos116_78 in116 sp78 11140.846016
Rwpos116_79 in116 sp79 3183.098862
Rwpos116_80 in116 sp80 11140.846016
Rwpos116_81 in116 sp81 3183.098862
Rwpos116_82 in116 sp82 3183.098862
Rwpos116_83 in116 sp83 11140.846016
Rwpos116_84 in116 sp84 11140.846016
Rwpos116_85 in116 sp85 3183.098862
Rwpos116_86 in116 sp86 11140.846016
Rwpos116_87 in116 sp87 3183.098862
Rwpos116_88 in116 sp88 3183.098862
Rwpos116_89 in116 sp89 3183.098862
Rwpos116_90 in116 sp90 3183.098862
Rwpos116_91 in116 sp91 3183.098862
Rwpos116_92 in116 sp92 11140.846016
Rwpos116_93 in116 sp93 3183.098862
Rwpos116_94 in116 sp94 11140.846016
Rwpos116_95 in116 sp95 3183.098862
Rwpos116_96 in116 sp96 3183.098862
Rwpos116_97 in116 sp97 11140.846016
Rwpos116_98 in116 sp98 11140.846016
Rwpos116_99 in116 sp99 3183.098862
Rwpos116_100 in116 sp100 3183.098862
Rwpos117_1 in117 sp1 3183.098862
Rwpos117_2 in117 sp2 11140.846016
Rwpos117_3 in117 sp3 11140.846016
Rwpos117_4 in117 sp4 11140.846016
Rwpos117_5 in117 sp5 11140.846016
Rwpos117_6 in117 sp6 11140.846016
Rwpos117_7 in117 sp7 3183.098862
Rwpos117_8 in117 sp8 3183.098862
Rwpos117_9 in117 sp9 11140.846016
Rwpos117_10 in117 sp10 11140.846016
Rwpos117_11 in117 sp11 3183.098862
Rwpos117_12 in117 sp12 11140.846016
Rwpos117_13 in117 sp13 3183.098862
Rwpos117_14 in117 sp14 11140.846016
Rwpos117_15 in117 sp15 3183.098862
Rwpos117_16 in117 sp16 11140.846016
Rwpos117_17 in117 sp17 3183.098862
Rwpos117_18 in117 sp18 11140.846016
Rwpos117_19 in117 sp19 3183.098862
Rwpos117_20 in117 sp20 11140.846016
Rwpos117_21 in117 sp21 3183.098862
Rwpos117_22 in117 sp22 3183.098862
Rwpos117_23 in117 sp23 3183.098862
Rwpos117_24 in117 sp24 11140.846016
Rwpos117_25 in117 sp25 11140.846016
Rwpos117_26 in117 sp26 11140.846016
Rwpos117_27 in117 sp27 3183.098862
Rwpos117_28 in117 sp28 3183.098862
Rwpos117_29 in117 sp29 3183.098862
Rwpos117_30 in117 sp30 3183.098862
Rwpos117_31 in117 sp31 11140.846016
Rwpos117_32 in117 sp32 11140.846016
Rwpos117_33 in117 sp33 11140.846016
Rwpos117_34 in117 sp34 3183.098862
Rwpos117_35 in117 sp35 3183.098862
Rwpos117_36 in117 sp36 3183.098862
Rwpos117_37 in117 sp37 3183.098862
Rwpos117_38 in117 sp38 3183.098862
Rwpos117_39 in117 sp39 11140.846016
Rwpos117_40 in117 sp40 3183.098862
Rwpos117_41 in117 sp41 3183.098862
Rwpos117_42 in117 sp42 11140.846016
Rwpos117_43 in117 sp43 3183.098862
Rwpos117_44 in117 sp44 11140.846016
Rwpos117_45 in117 sp45 11140.846016
Rwpos117_46 in117 sp46 11140.846016
Rwpos117_47 in117 sp47 3183.098862
Rwpos117_48 in117 sp48 11140.846016
Rwpos117_49 in117 sp49 11140.846016
Rwpos117_50 in117 sp50 3183.098862
Rwpos117_51 in117 sp51 3183.098862
Rwpos117_52 in117 sp52 11140.846016
Rwpos117_53 in117 sp53 3183.098862
Rwpos117_54 in117 sp54 3183.098862
Rwpos117_55 in117 sp55 11140.846016
Rwpos117_56 in117 sp56 3183.098862
Rwpos117_57 in117 sp57 3183.098862
Rwpos117_58 in117 sp58 11140.846016
Rwpos117_59 in117 sp59 11140.846016
Rwpos117_60 in117 sp60 11140.846016
Rwpos117_61 in117 sp61 3183.098862
Rwpos117_62 in117 sp62 3183.098862
Rwpos117_63 in117 sp63 3183.098862
Rwpos117_64 in117 sp64 11140.846016
Rwpos117_65 in117 sp65 11140.846016
Rwpos117_66 in117 sp66 11140.846016
Rwpos117_67 in117 sp67 3183.098862
Rwpos117_68 in117 sp68 11140.846016
Rwpos117_69 in117 sp69 11140.846016
Rwpos117_70 in117 sp70 3183.098862
Rwpos117_71 in117 sp71 3183.098862
Rwpos117_72 in117 sp72 11140.846016
Rwpos117_73 in117 sp73 3183.098862
Rwpos117_74 in117 sp74 11140.846016
Rwpos117_75 in117 sp75 3183.098862
Rwpos117_76 in117 sp76 11140.846016
Rwpos117_77 in117 sp77 11140.846016
Rwpos117_78 in117 sp78 11140.846016
Rwpos117_79 in117 sp79 3183.098862
Rwpos117_80 in117 sp80 11140.846016
Rwpos117_81 in117 sp81 3183.098862
Rwpos117_82 in117 sp82 3183.098862
Rwpos117_83 in117 sp83 11140.846016
Rwpos117_84 in117 sp84 11140.846016
Rwpos117_85 in117 sp85 3183.098862
Rwpos117_86 in117 sp86 3183.098862
Rwpos117_87 in117 sp87 3183.098862
Rwpos117_88 in117 sp88 3183.098862
Rwpos117_89 in117 sp89 11140.846016
Rwpos117_90 in117 sp90 3183.098862
Rwpos117_91 in117 sp91 11140.846016
Rwpos117_92 in117 sp92 11140.846016
Rwpos117_93 in117 sp93 11140.846016
Rwpos117_94 in117 sp94 3183.098862
Rwpos117_95 in117 sp95 11140.846016
Rwpos117_96 in117 sp96 11140.846016
Rwpos117_97 in117 sp97 3183.098862
Rwpos117_98 in117 sp98 3183.098862
Rwpos117_99 in117 sp99 11140.846016
Rwpos117_100 in117 sp100 11140.846016
Rwpos118_1 in118 sp1 3183.098862
Rwpos118_2 in118 sp2 3183.098862
Rwpos118_3 in118 sp3 11140.846016
Rwpos118_4 in118 sp4 3183.098862
Rwpos118_5 in118 sp5 11140.846016
Rwpos118_6 in118 sp6 3183.098862
Rwpos118_7 in118 sp7 11140.846016
Rwpos118_8 in118 sp8 11140.846016
Rwpos118_9 in118 sp9 11140.846016
Rwpos118_10 in118 sp10 3183.098862
Rwpos118_11 in118 sp11 3183.098862
Rwpos118_12 in118 sp12 11140.846016
Rwpos118_13 in118 sp13 11140.846016
Rwpos118_14 in118 sp14 3183.098862
Rwpos118_15 in118 sp15 3183.098862
Rwpos118_16 in118 sp16 3183.098862
Rwpos118_17 in118 sp17 11140.846016
Rwpos118_18 in118 sp18 3183.098862
Rwpos118_19 in118 sp19 3183.098862
Rwpos118_20 in118 sp20 3183.098862
Rwpos118_21 in118 sp21 3183.098862
Rwpos118_22 in118 sp22 11140.846016
Rwpos118_23 in118 sp23 11140.846016
Rwpos118_24 in118 sp24 11140.846016
Rwpos118_25 in118 sp25 11140.846016
Rwpos118_26 in118 sp26 11140.846016
Rwpos118_27 in118 sp27 3183.098862
Rwpos118_28 in118 sp28 3183.098862
Rwpos118_29 in118 sp29 3183.098862
Rwpos118_30 in118 sp30 3183.098862
Rwpos118_31 in118 sp31 3183.098862
Rwpos118_32 in118 sp32 11140.846016
Rwpos118_33 in118 sp33 3183.098862
Rwpos118_34 in118 sp34 11140.846016
Rwpos118_35 in118 sp35 11140.846016
Rwpos118_36 in118 sp36 3183.098862
Rwpos118_37 in118 sp37 3183.098862
Rwpos118_38 in118 sp38 3183.098862
Rwpos118_39 in118 sp39 11140.846016
Rwpos118_40 in118 sp40 3183.098862
Rwpos118_41 in118 sp41 3183.098862
Rwpos118_42 in118 sp42 11140.846016
Rwpos118_43 in118 sp43 11140.846016
Rwpos118_44 in118 sp44 3183.098862
Rwpos118_45 in118 sp45 3183.098862
Rwpos118_46 in118 sp46 3183.098862
Rwpos118_47 in118 sp47 3183.098862
Rwpos118_48 in118 sp48 11140.846016
Rwpos118_49 in118 sp49 11140.846016
Rwpos118_50 in118 sp50 3183.098862
Rwpos118_51 in118 sp51 11140.846016
Rwpos118_52 in118 sp52 3183.098862
Rwpos118_53 in118 sp53 3183.098862
Rwpos118_54 in118 sp54 11140.846016
Rwpos118_55 in118 sp55 11140.846016
Rwpos118_56 in118 sp56 3183.098862
Rwpos118_57 in118 sp57 11140.846016
Rwpos118_58 in118 sp58 3183.098862
Rwpos118_59 in118 sp59 11140.846016
Rwpos118_60 in118 sp60 11140.846016
Rwpos118_61 in118 sp61 11140.846016
Rwpos118_62 in118 sp62 11140.846016
Rwpos118_63 in118 sp63 11140.846016
Rwpos118_64 in118 sp64 11140.846016
Rwpos118_65 in118 sp65 3183.098862
Rwpos118_66 in118 sp66 11140.846016
Rwpos118_67 in118 sp67 3183.098862
Rwpos118_68 in118 sp68 11140.846016
Rwpos118_69 in118 sp69 11140.846016
Rwpos118_70 in118 sp70 11140.846016
Rwpos118_71 in118 sp71 3183.098862
Rwpos118_72 in118 sp72 3183.098862
Rwpos118_73 in118 sp73 3183.098862
Rwpos118_74 in118 sp74 3183.098862
Rwpos118_75 in118 sp75 3183.098862
Rwpos118_76 in118 sp76 11140.846016
Rwpos118_77 in118 sp77 11140.846016
Rwpos118_78 in118 sp78 11140.846016
Rwpos118_79 in118 sp79 3183.098862
Rwpos118_80 in118 sp80 11140.846016
Rwpos118_81 in118 sp81 3183.098862
Rwpos118_82 in118 sp82 3183.098862
Rwpos118_83 in118 sp83 3183.098862
Rwpos118_84 in118 sp84 11140.846016
Rwpos118_85 in118 sp85 11140.846016
Rwpos118_86 in118 sp86 11140.846016
Rwpos118_87 in118 sp87 11140.846016
Rwpos118_88 in118 sp88 3183.098862
Rwpos118_89 in118 sp89 11140.846016
Rwpos118_90 in118 sp90 3183.098862
Rwpos118_91 in118 sp91 3183.098862
Rwpos118_92 in118 sp92 11140.846016
Rwpos118_93 in118 sp93 3183.098862
Rwpos118_94 in118 sp94 3183.098862
Rwpos118_95 in118 sp95 11140.846016
Rwpos118_96 in118 sp96 3183.098862
Rwpos118_97 in118 sp97 11140.846016
Rwpos118_98 in118 sp98 11140.846016
Rwpos118_99 in118 sp99 11140.846016
Rwpos118_100 in118 sp100 11140.846016
Rwpos119_1 in119 sp1 3183.098862
Rwpos119_2 in119 sp2 3183.098862
Rwpos119_3 in119 sp3 11140.846016
Rwpos119_4 in119 sp4 11140.846016
Rwpos119_5 in119 sp5 3183.098862
Rwpos119_6 in119 sp6 11140.846016
Rwpos119_7 in119 sp7 11140.846016
Rwpos119_8 in119 sp8 3183.098862
Rwpos119_9 in119 sp9 11140.846016
Rwpos119_10 in119 sp10 3183.098862
Rwpos119_11 in119 sp11 11140.846016
Rwpos119_12 in119 sp12 3183.098862
Rwpos119_13 in119 sp13 11140.846016
Rwpos119_14 in119 sp14 3183.098862
Rwpos119_15 in119 sp15 3183.098862
Rwpos119_16 in119 sp16 3183.098862
Rwpos119_17 in119 sp17 3183.098862
Rwpos119_18 in119 sp18 11140.846016
Rwpos119_19 in119 sp19 11140.846016
Rwpos119_20 in119 sp20 3183.098862
Rwpos119_21 in119 sp21 3183.098862
Rwpos119_22 in119 sp22 11140.846016
Rwpos119_23 in119 sp23 11140.846016
Rwpos119_24 in119 sp24 3183.098862
Rwpos119_25 in119 sp25 11140.846016
Rwpos119_26 in119 sp26 3183.098862
Rwpos119_27 in119 sp27 3183.098862
Rwpos119_28 in119 sp28 11140.846016
Rwpos119_29 in119 sp29 3183.098862
Rwpos119_30 in119 sp30 3183.098862
Rwpos119_31 in119 sp31 11140.846016
Rwpos119_32 in119 sp32 3183.098862
Rwpos119_33 in119 sp33 3183.098862
Rwpos119_34 in119 sp34 3183.098862
Rwpos119_35 in119 sp35 3183.098862
Rwpos119_36 in119 sp36 3183.098862
Rwpos119_37 in119 sp37 11140.846016
Rwpos119_38 in119 sp38 3183.098862
Rwpos119_39 in119 sp39 3183.098862
Rwpos119_40 in119 sp40 3183.098862
Rwpos119_41 in119 sp41 11140.846016
Rwpos119_42 in119 sp42 3183.098862
Rwpos119_43 in119 sp43 11140.846016
Rwpos119_44 in119 sp44 3183.098862
Rwpos119_45 in119 sp45 11140.846016
Rwpos119_46 in119 sp46 3183.098862
Rwpos119_47 in119 sp47 3183.098862
Rwpos119_48 in119 sp48 3183.098862
Rwpos119_49 in119 sp49 3183.098862
Rwpos119_50 in119 sp50 3183.098862
Rwpos119_51 in119 sp51 3183.098862
Rwpos119_52 in119 sp52 3183.098862
Rwpos119_53 in119 sp53 11140.846016
Rwpos119_54 in119 sp54 3183.098862
Rwpos119_55 in119 sp55 3183.098862
Rwpos119_56 in119 sp56 3183.098862
Rwpos119_57 in119 sp57 11140.846016
Rwpos119_58 in119 sp58 3183.098862
Rwpos119_59 in119 sp59 11140.846016
Rwpos119_60 in119 sp60 11140.846016
Rwpos119_61 in119 sp61 11140.846016
Rwpos119_62 in119 sp62 3183.098862
Rwpos119_63 in119 sp63 3183.098862
Rwpos119_64 in119 sp64 11140.846016
Rwpos119_65 in119 sp65 11140.846016
Rwpos119_66 in119 sp66 3183.098862
Rwpos119_67 in119 sp67 3183.098862
Rwpos119_68 in119 sp68 3183.098862
Rwpos119_69 in119 sp69 3183.098862
Rwpos119_70 in119 sp70 3183.098862
Rwpos119_71 in119 sp71 11140.846016
Rwpos119_72 in119 sp72 11140.846016
Rwpos119_73 in119 sp73 11140.846016
Rwpos119_74 in119 sp74 3183.098862
Rwpos119_75 in119 sp75 11140.846016
Rwpos119_76 in119 sp76 11140.846016
Rwpos119_77 in119 sp77 11140.846016
Rwpos119_78 in119 sp78 11140.846016
Rwpos119_79 in119 sp79 3183.098862
Rwpos119_80 in119 sp80 11140.846016
Rwpos119_81 in119 sp81 11140.846016
Rwpos119_82 in119 sp82 3183.098862
Rwpos119_83 in119 sp83 11140.846016
Rwpos119_84 in119 sp84 11140.846016
Rwpos119_85 in119 sp85 3183.098862
Rwpos119_86 in119 sp86 11140.846016
Rwpos119_87 in119 sp87 3183.098862
Rwpos119_88 in119 sp88 3183.098862
Rwpos119_89 in119 sp89 11140.846016
Rwpos119_90 in119 sp90 3183.098862
Rwpos119_91 in119 sp91 11140.846016
Rwpos119_92 in119 sp92 11140.846016
Rwpos119_93 in119 sp93 11140.846016
Rwpos119_94 in119 sp94 3183.098862
Rwpos119_95 in119 sp95 3183.098862
Rwpos119_96 in119 sp96 11140.846016
Rwpos119_97 in119 sp97 11140.846016
Rwpos119_98 in119 sp98 3183.098862
Rwpos119_99 in119 sp99 3183.098862
Rwpos119_100 in119 sp100 3183.098862
Rwpos120_1 in120 sp1 3183.098862
Rwpos120_2 in120 sp2 3183.098862
Rwpos120_3 in120 sp3 11140.846016
Rwpos120_4 in120 sp4 3183.098862
Rwpos120_5 in120 sp5 11140.846016
Rwpos120_6 in120 sp6 3183.098862
Rwpos120_7 in120 sp7 11140.846016
Rwpos120_8 in120 sp8 3183.098862
Rwpos120_9 in120 sp9 3183.098862
Rwpos120_10 in120 sp10 3183.098862
Rwpos120_11 in120 sp11 3183.098862
Rwpos120_12 in120 sp12 11140.846016
Rwpos120_13 in120 sp13 11140.846016
Rwpos120_14 in120 sp14 3183.098862
Rwpos120_15 in120 sp15 3183.098862
Rwpos120_16 in120 sp16 3183.098862
Rwpos120_17 in120 sp17 3183.098862
Rwpos120_18 in120 sp18 3183.098862
Rwpos120_19 in120 sp19 11140.846016
Rwpos120_20 in120 sp20 3183.098862
Rwpos120_21 in120 sp21 11140.846016
Rwpos120_22 in120 sp22 3183.098862
Rwpos120_23 in120 sp23 11140.846016
Rwpos120_24 in120 sp24 11140.846016
Rwpos120_25 in120 sp25 11140.846016
Rwpos120_26 in120 sp26 3183.098862
Rwpos120_27 in120 sp27 3183.098862
Rwpos120_28 in120 sp28 11140.846016
Rwpos120_29 in120 sp29 3183.098862
Rwpos120_30 in120 sp30 3183.098862
Rwpos120_31 in120 sp31 3183.098862
Rwpos120_32 in120 sp32 3183.098862
Rwpos120_33 in120 sp33 3183.098862
Rwpos120_34 in120 sp34 3183.098862
Rwpos120_35 in120 sp35 11140.846016
Rwpos120_36 in120 sp36 3183.098862
Rwpos120_37 in120 sp37 11140.846016
Rwpos120_38 in120 sp38 3183.098862
Rwpos120_39 in120 sp39 11140.846016
Rwpos120_40 in120 sp40 11140.846016
Rwpos120_41 in120 sp41 11140.846016
Rwpos120_42 in120 sp42 11140.846016
Rwpos120_43 in120 sp43 3183.098862
Rwpos120_44 in120 sp44 3183.098862
Rwpos120_45 in120 sp45 3183.098862
Rwpos120_46 in120 sp46 3183.098862
Rwpos120_47 in120 sp47 3183.098862
Rwpos120_48 in120 sp48 3183.098862
Rwpos120_49 in120 sp49 3183.098862
Rwpos120_50 in120 sp50 3183.098862
Rwpos120_51 in120 sp51 11140.846016
Rwpos120_52 in120 sp52 11140.846016
Rwpos120_53 in120 sp53 3183.098862
Rwpos120_54 in120 sp54 3183.098862
Rwpos120_55 in120 sp55 3183.098862
Rwpos120_56 in120 sp56 3183.098862
Rwpos120_57 in120 sp57 11140.846016
Rwpos120_58 in120 sp58 3183.098862
Rwpos120_59 in120 sp59 11140.846016
Rwpos120_60 in120 sp60 3183.098862
Rwpos120_61 in120 sp61 3183.098862
Rwpos120_62 in120 sp62 11140.846016
Rwpos120_63 in120 sp63 3183.098862
Rwpos120_64 in120 sp64 3183.098862
Rwpos120_65 in120 sp65 3183.098862
Rwpos120_66 in120 sp66 11140.846016
Rwpos120_67 in120 sp67 3183.098862
Rwpos120_68 in120 sp68 3183.098862
Rwpos120_69 in120 sp69 3183.098862
Rwpos120_70 in120 sp70 3183.098862
Rwpos120_71 in120 sp71 11140.846016
Rwpos120_72 in120 sp72 11140.846016
Rwpos120_73 in120 sp73 11140.846016
Rwpos120_74 in120 sp74 11140.846016
Rwpos120_75 in120 sp75 11140.846016
Rwpos120_76 in120 sp76 3183.098862
Rwpos120_77 in120 sp77 11140.846016
Rwpos120_78 in120 sp78 3183.098862
Rwpos120_79 in120 sp79 11140.846016
Rwpos120_80 in120 sp80 11140.846016
Rwpos120_81 in120 sp81 11140.846016
Rwpos120_82 in120 sp82 3183.098862
Rwpos120_83 in120 sp83 11140.846016
Rwpos120_84 in120 sp84 11140.846016
Rwpos120_85 in120 sp85 3183.098862
Rwpos120_86 in120 sp86 11140.846016
Rwpos120_87 in120 sp87 3183.098862
Rwpos120_88 in120 sp88 11140.846016
Rwpos120_89 in120 sp89 11140.846016
Rwpos120_90 in120 sp90 3183.098862
Rwpos120_91 in120 sp91 3183.098862
Rwpos120_92 in120 sp92 11140.846016
Rwpos120_93 in120 sp93 3183.098862
Rwpos120_94 in120 sp94 3183.098862
Rwpos120_95 in120 sp95 11140.846016
Rwpos120_96 in120 sp96 3183.098862
Rwpos120_97 in120 sp97 3183.098862
Rwpos120_98 in120 sp98 11140.846016
Rwpos120_99 in120 sp99 11140.846016
Rwpos120_100 in120 sp100 3183.098862
Rwpos121_1 in121 sp1 11140.846016
Rwpos121_2 in121 sp2 11140.846016
Rwpos121_3 in121 sp3 3183.098862
Rwpos121_4 in121 sp4 3183.098862
Rwpos121_5 in121 sp5 11140.846016
Rwpos121_6 in121 sp6 3183.098862
Rwpos121_7 in121 sp7 11140.846016
Rwpos121_8 in121 sp8 3183.098862
Rwpos121_9 in121 sp9 3183.098862
Rwpos121_10 in121 sp10 3183.098862
Rwpos121_11 in121 sp11 3183.098862
Rwpos121_12 in121 sp12 11140.846016
Rwpos121_13 in121 sp13 3183.098862
Rwpos121_14 in121 sp14 11140.846016
Rwpos121_15 in121 sp15 3183.098862
Rwpos121_16 in121 sp16 11140.846016
Rwpos121_17 in121 sp17 11140.846016
Rwpos121_18 in121 sp18 11140.846016
Rwpos121_19 in121 sp19 3183.098862
Rwpos121_20 in121 sp20 3183.098862
Rwpos121_21 in121 sp21 3183.098862
Rwpos121_22 in121 sp22 3183.098862
Rwpos121_23 in121 sp23 11140.846016
Rwpos121_24 in121 sp24 3183.098862
Rwpos121_25 in121 sp25 11140.846016
Rwpos121_26 in121 sp26 11140.846016
Rwpos121_27 in121 sp27 11140.846016
Rwpos121_28 in121 sp28 11140.846016
Rwpos121_29 in121 sp29 11140.846016
Rwpos121_30 in121 sp30 11140.846016
Rwpos121_31 in121 sp31 3183.098862
Rwpos121_32 in121 sp32 11140.846016
Rwpos121_33 in121 sp33 3183.098862
Rwpos121_34 in121 sp34 11140.846016
Rwpos121_35 in121 sp35 3183.098862
Rwpos121_36 in121 sp36 3183.098862
Rwpos121_37 in121 sp37 3183.098862
Rwpos121_38 in121 sp38 11140.846016
Rwpos121_39 in121 sp39 3183.098862
Rwpos121_40 in121 sp40 3183.098862
Rwpos121_41 in121 sp41 3183.098862
Rwpos121_42 in121 sp42 11140.846016
Rwpos121_43 in121 sp43 3183.098862
Rwpos121_44 in121 sp44 11140.846016
Rwpos121_45 in121 sp45 11140.846016
Rwpos121_46 in121 sp46 11140.846016
Rwpos121_47 in121 sp47 11140.846016
Rwpos121_48 in121 sp48 11140.846016
Rwpos121_49 in121 sp49 3183.098862
Rwpos121_50 in121 sp50 11140.846016
Rwpos121_51 in121 sp51 11140.846016
Rwpos121_52 in121 sp52 3183.098862
Rwpos121_53 in121 sp53 11140.846016
Rwpos121_54 in121 sp54 3183.098862
Rwpos121_55 in121 sp55 11140.846016
Rwpos121_56 in121 sp56 3183.098862
Rwpos121_57 in121 sp57 11140.846016
Rwpos121_58 in121 sp58 3183.098862
Rwpos121_59 in121 sp59 11140.846016
Rwpos121_60 in121 sp60 3183.098862
Rwpos121_61 in121 sp61 11140.846016
Rwpos121_62 in121 sp62 11140.846016
Rwpos121_63 in121 sp63 11140.846016
Rwpos121_64 in121 sp64 11140.846016
Rwpos121_65 in121 sp65 3183.098862
Rwpos121_66 in121 sp66 11140.846016
Rwpos121_67 in121 sp67 3183.098862
Rwpos121_68 in121 sp68 3183.098862
Rwpos121_69 in121 sp69 11140.846016
Rwpos121_70 in121 sp70 3183.098862
Rwpos121_71 in121 sp71 3183.098862
Rwpos121_72 in121 sp72 3183.098862
Rwpos121_73 in121 sp73 3183.098862
Rwpos121_74 in121 sp74 3183.098862
Rwpos121_75 in121 sp75 3183.098862
Rwpos121_76 in121 sp76 11140.846016
Rwpos121_77 in121 sp77 11140.846016
Rwpos121_78 in121 sp78 3183.098862
Rwpos121_79 in121 sp79 3183.098862
Rwpos121_80 in121 sp80 11140.846016
Rwpos121_81 in121 sp81 11140.846016
Rwpos121_82 in121 sp82 11140.846016
Rwpos121_83 in121 sp83 3183.098862
Rwpos121_84 in121 sp84 3183.098862
Rwpos121_85 in121 sp85 3183.098862
Rwpos121_86 in121 sp86 11140.846016
Rwpos121_87 in121 sp87 11140.846016
Rwpos121_88 in121 sp88 11140.846016
Rwpos121_89 in121 sp89 3183.098862
Rwpos121_90 in121 sp90 3183.098862
Rwpos121_91 in121 sp91 3183.098862
Rwpos121_92 in121 sp92 3183.098862
Rwpos121_93 in121 sp93 3183.098862
Rwpos121_94 in121 sp94 11140.846016
Rwpos121_95 in121 sp95 3183.098862
Rwpos121_96 in121 sp96 3183.098862
Rwpos121_97 in121 sp97 3183.098862
Rwpos121_98 in121 sp98 3183.098862
Rwpos121_99 in121 sp99 3183.098862
Rwpos121_100 in121 sp100 11140.846016
Rwpos122_1 in122 sp1 3183.098862
Rwpos122_2 in122 sp2 11140.846016
Rwpos122_3 in122 sp3 11140.846016
Rwpos122_4 in122 sp4 3183.098862
Rwpos122_5 in122 sp5 3183.098862
Rwpos122_6 in122 sp6 11140.846016
Rwpos122_7 in122 sp7 11140.846016
Rwpos122_8 in122 sp8 3183.098862
Rwpos122_9 in122 sp9 3183.098862
Rwpos122_10 in122 sp10 11140.846016
Rwpos122_11 in122 sp11 11140.846016
Rwpos122_12 in122 sp12 11140.846016
Rwpos122_13 in122 sp13 3183.098862
Rwpos122_14 in122 sp14 11140.846016
Rwpos122_15 in122 sp15 3183.098862
Rwpos122_16 in122 sp16 11140.846016
Rwpos122_17 in122 sp17 3183.098862
Rwpos122_18 in122 sp18 11140.846016
Rwpos122_19 in122 sp19 3183.098862
Rwpos122_20 in122 sp20 3183.098862
Rwpos122_21 in122 sp21 11140.846016
Rwpos122_22 in122 sp22 3183.098862
Rwpos122_23 in122 sp23 11140.846016
Rwpos122_24 in122 sp24 11140.846016
Rwpos122_25 in122 sp25 11140.846016
Rwpos122_26 in122 sp26 11140.846016
Rwpos122_27 in122 sp27 3183.098862
Rwpos122_28 in122 sp28 3183.098862
Rwpos122_29 in122 sp29 11140.846016
Rwpos122_30 in122 sp30 11140.846016
Rwpos122_31 in122 sp31 11140.846016
Rwpos122_32 in122 sp32 3183.098862
Rwpos122_33 in122 sp33 3183.098862
Rwpos122_34 in122 sp34 11140.846016
Rwpos122_35 in122 sp35 3183.098862
Rwpos122_36 in122 sp36 3183.098862
Rwpos122_37 in122 sp37 3183.098862
Rwpos122_38 in122 sp38 11140.846016
Rwpos122_39 in122 sp39 11140.846016
Rwpos122_40 in122 sp40 3183.098862
Rwpos122_41 in122 sp41 3183.098862
Rwpos122_42 in122 sp42 11140.846016
Rwpos122_43 in122 sp43 3183.098862
Rwpos122_44 in122 sp44 3183.098862
Rwpos122_45 in122 sp45 11140.846016
Rwpos122_46 in122 sp46 11140.846016
Rwpos122_47 in122 sp47 11140.846016
Rwpos122_48 in122 sp48 3183.098862
Rwpos122_49 in122 sp49 3183.098862
Rwpos122_50 in122 sp50 3183.098862
Rwpos122_51 in122 sp51 11140.846016
Rwpos122_52 in122 sp52 3183.098862
Rwpos122_53 in122 sp53 11140.846016
Rwpos122_54 in122 sp54 11140.846016
Rwpos122_55 in122 sp55 3183.098862
Rwpos122_56 in122 sp56 3183.098862
Rwpos122_57 in122 sp57 11140.846016
Rwpos122_58 in122 sp58 11140.846016
Rwpos122_59 in122 sp59 3183.098862
Rwpos122_60 in122 sp60 11140.846016
Rwpos122_61 in122 sp61 3183.098862
Rwpos122_62 in122 sp62 11140.846016
Rwpos122_63 in122 sp63 3183.098862
Rwpos122_64 in122 sp64 11140.846016
Rwpos122_65 in122 sp65 11140.846016
Rwpos122_66 in122 sp66 3183.098862
Rwpos122_67 in122 sp67 3183.098862
Rwpos122_68 in122 sp68 11140.846016
Rwpos122_69 in122 sp69 11140.846016
Rwpos122_70 in122 sp70 3183.098862
Rwpos122_71 in122 sp71 11140.846016
Rwpos122_72 in122 sp72 3183.098862
Rwpos122_73 in122 sp73 3183.098862
Rwpos122_74 in122 sp74 11140.846016
Rwpos122_75 in122 sp75 3183.098862
Rwpos122_76 in122 sp76 3183.098862
Rwpos122_77 in122 sp77 11140.846016
Rwpos122_78 in122 sp78 3183.098862
Rwpos122_79 in122 sp79 3183.098862
Rwpos122_80 in122 sp80 11140.846016
Rwpos122_81 in122 sp81 3183.098862
Rwpos122_82 in122 sp82 3183.098862
Rwpos122_83 in122 sp83 11140.846016
Rwpos122_84 in122 sp84 3183.098862
Rwpos122_85 in122 sp85 3183.098862
Rwpos122_86 in122 sp86 11140.846016
Rwpos122_87 in122 sp87 3183.098862
Rwpos122_88 in122 sp88 11140.846016
Rwpos122_89 in122 sp89 11140.846016
Rwpos122_90 in122 sp90 11140.846016
Rwpos122_91 in122 sp91 3183.098862
Rwpos122_92 in122 sp92 3183.098862
Rwpos122_93 in122 sp93 3183.098862
Rwpos122_94 in122 sp94 3183.098862
Rwpos122_95 in122 sp95 11140.846016
Rwpos122_96 in122 sp96 11140.846016
Rwpos122_97 in122 sp97 3183.098862
Rwpos122_98 in122 sp98 11140.846016
Rwpos122_99 in122 sp99 11140.846016
Rwpos122_100 in122 sp100 11140.846016
Rwpos123_1 in123 sp1 11140.846016
Rwpos123_2 in123 sp2 11140.846016
Rwpos123_3 in123 sp3 11140.846016
Rwpos123_4 in123 sp4 11140.846016
Rwpos123_5 in123 sp5 11140.846016
Rwpos123_6 in123 sp6 3183.098862
Rwpos123_7 in123 sp7 3183.098862
Rwpos123_8 in123 sp8 11140.846016
Rwpos123_9 in123 sp9 11140.846016
Rwpos123_10 in123 sp10 3183.098862
Rwpos123_11 in123 sp11 11140.846016
Rwpos123_12 in123 sp12 11140.846016
Rwpos123_13 in123 sp13 11140.846016
Rwpos123_14 in123 sp14 3183.098862
Rwpos123_15 in123 sp15 3183.098862
Rwpos123_16 in123 sp16 11140.846016
Rwpos123_17 in123 sp17 11140.846016
Rwpos123_18 in123 sp18 11140.846016
Rwpos123_19 in123 sp19 11140.846016
Rwpos123_20 in123 sp20 11140.846016
Rwpos123_21 in123 sp21 11140.846016
Rwpos123_22 in123 sp22 11140.846016
Rwpos123_23 in123 sp23 11140.846016
Rwpos123_24 in123 sp24 11140.846016
Rwpos123_25 in123 sp25 11140.846016
Rwpos123_26 in123 sp26 3183.098862
Rwpos123_27 in123 sp27 3183.098862
Rwpos123_28 in123 sp28 3183.098862
Rwpos123_29 in123 sp29 3183.098862
Rwpos123_30 in123 sp30 3183.098862
Rwpos123_31 in123 sp31 11140.846016
Rwpos123_32 in123 sp32 3183.098862
Rwpos123_33 in123 sp33 3183.098862
Rwpos123_34 in123 sp34 3183.098862
Rwpos123_35 in123 sp35 3183.098862
Rwpos123_36 in123 sp36 3183.098862
Rwpos123_37 in123 sp37 3183.098862
Rwpos123_38 in123 sp38 11140.846016
Rwpos123_39 in123 sp39 3183.098862
Rwpos123_40 in123 sp40 11140.846016
Rwpos123_41 in123 sp41 3183.098862
Rwpos123_42 in123 sp42 3183.098862
Rwpos123_43 in123 sp43 3183.098862
Rwpos123_44 in123 sp44 3183.098862
Rwpos123_45 in123 sp45 11140.846016
Rwpos123_46 in123 sp46 3183.098862
Rwpos123_47 in123 sp47 11140.846016
Rwpos123_48 in123 sp48 3183.098862
Rwpos123_49 in123 sp49 11140.846016
Rwpos123_50 in123 sp50 11140.846016
Rwpos123_51 in123 sp51 11140.846016
Rwpos123_52 in123 sp52 11140.846016
Rwpos123_53 in123 sp53 3183.098862
Rwpos123_54 in123 sp54 11140.846016
Rwpos123_55 in123 sp55 11140.846016
Rwpos123_56 in123 sp56 3183.098862
Rwpos123_57 in123 sp57 3183.098862
Rwpos123_58 in123 sp58 11140.846016
Rwpos123_59 in123 sp59 11140.846016
Rwpos123_60 in123 sp60 11140.846016
Rwpos123_61 in123 sp61 3183.098862
Rwpos123_62 in123 sp62 3183.098862
Rwpos123_63 in123 sp63 11140.846016
Rwpos123_64 in123 sp64 3183.098862
Rwpos123_65 in123 sp65 11140.846016
Rwpos123_66 in123 sp66 11140.846016
Rwpos123_67 in123 sp67 3183.098862
Rwpos123_68 in123 sp68 11140.846016
Rwpos123_69 in123 sp69 11140.846016
Rwpos123_70 in123 sp70 3183.098862
Rwpos123_71 in123 sp71 3183.098862
Rwpos123_72 in123 sp72 11140.846016
Rwpos123_73 in123 sp73 11140.846016
Rwpos123_74 in123 sp74 11140.846016
Rwpos123_75 in123 sp75 3183.098862
Rwpos123_76 in123 sp76 3183.098862
Rwpos123_77 in123 sp77 3183.098862
Rwpos123_78 in123 sp78 11140.846016
Rwpos123_79 in123 sp79 3183.098862
Rwpos123_80 in123 sp80 3183.098862
Rwpos123_81 in123 sp81 11140.846016
Rwpos123_82 in123 sp82 11140.846016
Rwpos123_83 in123 sp83 11140.846016
Rwpos123_84 in123 sp84 11140.846016
Rwpos123_85 in123 sp85 3183.098862
Rwpos123_86 in123 sp86 11140.846016
Rwpos123_87 in123 sp87 3183.098862
Rwpos123_88 in123 sp88 3183.098862
Rwpos123_89 in123 sp89 3183.098862
Rwpos123_90 in123 sp90 11140.846016
Rwpos123_91 in123 sp91 3183.098862
Rwpos123_92 in123 sp92 11140.846016
Rwpos123_93 in123 sp93 11140.846016
Rwpos123_94 in123 sp94 11140.846016
Rwpos123_95 in123 sp95 3183.098862
Rwpos123_96 in123 sp96 11140.846016
Rwpos123_97 in123 sp97 11140.846016
Rwpos123_98 in123 sp98 11140.846016
Rwpos123_99 in123 sp99 3183.098862
Rwpos123_100 in123 sp100 3183.098862
Rwpos124_1 in124 sp1 11140.846016
Rwpos124_2 in124 sp2 11140.846016
Rwpos124_3 in124 sp3 11140.846016
Rwpos124_4 in124 sp4 11140.846016
Rwpos124_5 in124 sp5 3183.098862
Rwpos124_6 in124 sp6 3183.098862
Rwpos124_7 in124 sp7 11140.846016
Rwpos124_8 in124 sp8 3183.098862
Rwpos124_9 in124 sp9 11140.846016
Rwpos124_10 in124 sp10 11140.846016
Rwpos124_11 in124 sp11 11140.846016
Rwpos124_12 in124 sp12 11140.846016
Rwpos124_13 in124 sp13 11140.846016
Rwpos124_14 in124 sp14 3183.098862
Rwpos124_15 in124 sp15 11140.846016
Rwpos124_16 in124 sp16 3183.098862
Rwpos124_17 in124 sp17 3183.098862
Rwpos124_18 in124 sp18 11140.846016
Rwpos124_19 in124 sp19 3183.098862
Rwpos124_20 in124 sp20 11140.846016
Rwpos124_21 in124 sp21 3183.098862
Rwpos124_22 in124 sp22 3183.098862
Rwpos124_23 in124 sp23 11140.846016
Rwpos124_24 in124 sp24 3183.098862
Rwpos124_25 in124 sp25 3183.098862
Rwpos124_26 in124 sp26 3183.098862
Rwpos124_27 in124 sp27 11140.846016
Rwpos124_28 in124 sp28 3183.098862
Rwpos124_29 in124 sp29 3183.098862
Rwpos124_30 in124 sp30 3183.098862
Rwpos124_31 in124 sp31 3183.098862
Rwpos124_32 in124 sp32 11140.846016
Rwpos124_33 in124 sp33 11140.846016
Rwpos124_34 in124 sp34 3183.098862
Rwpos124_35 in124 sp35 11140.846016
Rwpos124_36 in124 sp36 3183.098862
Rwpos124_37 in124 sp37 11140.846016
Rwpos124_38 in124 sp38 3183.098862
Rwpos124_39 in124 sp39 11140.846016
Rwpos124_40 in124 sp40 11140.846016
Rwpos124_41 in124 sp41 11140.846016
Rwpos124_42 in124 sp42 11140.846016
Rwpos124_43 in124 sp43 11140.846016
Rwpos124_44 in124 sp44 11140.846016
Rwpos124_45 in124 sp45 11140.846016
Rwpos124_46 in124 sp46 11140.846016
Rwpos124_47 in124 sp47 11140.846016
Rwpos124_48 in124 sp48 11140.846016
Rwpos124_49 in124 sp49 11140.846016
Rwpos124_50 in124 sp50 3183.098862
Rwpos124_51 in124 sp51 11140.846016
Rwpos124_52 in124 sp52 11140.846016
Rwpos124_53 in124 sp53 3183.098862
Rwpos124_54 in124 sp54 3183.098862
Rwpos124_55 in124 sp55 3183.098862
Rwpos124_56 in124 sp56 11140.846016
Rwpos124_57 in124 sp57 3183.098862
Rwpos124_58 in124 sp58 3183.098862
Rwpos124_59 in124 sp59 11140.846016
Rwpos124_60 in124 sp60 3183.098862
Rwpos124_61 in124 sp61 11140.846016
Rwpos124_62 in124 sp62 11140.846016
Rwpos124_63 in124 sp63 11140.846016
Rwpos124_64 in124 sp64 11140.846016
Rwpos124_65 in124 sp65 11140.846016
Rwpos124_66 in124 sp66 3183.098862
Rwpos124_67 in124 sp67 3183.098862
Rwpos124_68 in124 sp68 11140.846016
Rwpos124_69 in124 sp69 11140.846016
Rwpos124_70 in124 sp70 11140.846016
Rwpos124_71 in124 sp71 11140.846016
Rwpos124_72 in124 sp72 11140.846016
Rwpos124_73 in124 sp73 3183.098862
Rwpos124_74 in124 sp74 3183.098862
Rwpos124_75 in124 sp75 11140.846016
Rwpos124_76 in124 sp76 11140.846016
Rwpos124_77 in124 sp77 11140.846016
Rwpos124_78 in124 sp78 11140.846016
Rwpos124_79 in124 sp79 11140.846016
Rwpos124_80 in124 sp80 3183.098862
Rwpos124_81 in124 sp81 11140.846016
Rwpos124_82 in124 sp82 11140.846016
Rwpos124_83 in124 sp83 3183.098862
Rwpos124_84 in124 sp84 3183.098862
Rwpos124_85 in124 sp85 11140.846016
Rwpos124_86 in124 sp86 11140.846016
Rwpos124_87 in124 sp87 11140.846016
Rwpos124_88 in124 sp88 3183.098862
Rwpos124_89 in124 sp89 3183.098862
Rwpos124_90 in124 sp90 11140.846016
Rwpos124_91 in124 sp91 11140.846016
Rwpos124_92 in124 sp92 11140.846016
Rwpos124_93 in124 sp93 11140.846016
Rwpos124_94 in124 sp94 3183.098862
Rwpos124_95 in124 sp95 11140.846016
Rwpos124_96 in124 sp96 11140.846016
Rwpos124_97 in124 sp97 3183.098862
Rwpos124_98 in124 sp98 11140.846016
Rwpos124_99 in124 sp99 11140.846016
Rwpos124_100 in124 sp100 3183.098862
Rwpos125_1 in125 sp1 11140.846016
Rwpos125_2 in125 sp2 3183.098862
Rwpos125_3 in125 sp3 11140.846016
Rwpos125_4 in125 sp4 11140.846016
Rwpos125_5 in125 sp5 3183.098862
Rwpos125_6 in125 sp6 11140.846016
Rwpos125_7 in125 sp7 3183.098862
Rwpos125_8 in125 sp8 3183.098862
Rwpos125_9 in125 sp9 3183.098862
Rwpos125_10 in125 sp10 3183.098862
Rwpos125_11 in125 sp11 11140.846016
Rwpos125_12 in125 sp12 3183.098862
Rwpos125_13 in125 sp13 11140.846016
Rwpos125_14 in125 sp14 3183.098862
Rwpos125_15 in125 sp15 3183.098862
Rwpos125_16 in125 sp16 11140.846016
Rwpos125_17 in125 sp17 11140.846016
Rwpos125_18 in125 sp18 11140.846016
Rwpos125_19 in125 sp19 3183.098862
Rwpos125_20 in125 sp20 3183.098862
Rwpos125_21 in125 sp21 3183.098862
Rwpos125_22 in125 sp22 11140.846016
Rwpos125_23 in125 sp23 11140.846016
Rwpos125_24 in125 sp24 3183.098862
Rwpos125_25 in125 sp25 11140.846016
Rwpos125_26 in125 sp26 11140.846016
Rwpos125_27 in125 sp27 3183.098862
Rwpos125_28 in125 sp28 3183.098862
Rwpos125_29 in125 sp29 11140.846016
Rwpos125_30 in125 sp30 11140.846016
Rwpos125_31 in125 sp31 11140.846016
Rwpos125_32 in125 sp32 11140.846016
Rwpos125_33 in125 sp33 11140.846016
Rwpos125_34 in125 sp34 11140.846016
Rwpos125_35 in125 sp35 11140.846016
Rwpos125_36 in125 sp36 3183.098862
Rwpos125_37 in125 sp37 11140.846016
Rwpos125_38 in125 sp38 3183.098862
Rwpos125_39 in125 sp39 11140.846016
Rwpos125_40 in125 sp40 3183.098862
Rwpos125_41 in125 sp41 11140.846016
Rwpos125_42 in125 sp42 11140.846016
Rwpos125_43 in125 sp43 3183.098862
Rwpos125_44 in125 sp44 11140.846016
Rwpos125_45 in125 sp45 11140.846016
Rwpos125_46 in125 sp46 11140.846016
Rwpos125_47 in125 sp47 11140.846016
Rwpos125_48 in125 sp48 11140.846016
Rwpos125_49 in125 sp49 11140.846016
Rwpos125_50 in125 sp50 3183.098862
Rwpos125_51 in125 sp51 11140.846016
Rwpos125_52 in125 sp52 11140.846016
Rwpos125_53 in125 sp53 11140.846016
Rwpos125_54 in125 sp54 3183.098862
Rwpos125_55 in125 sp55 3183.098862
Rwpos125_56 in125 sp56 3183.098862
Rwpos125_57 in125 sp57 3183.098862
Rwpos125_58 in125 sp58 11140.846016
Rwpos125_59 in125 sp59 3183.098862
Rwpos125_60 in125 sp60 11140.846016
Rwpos125_61 in125 sp61 3183.098862
Rwpos125_62 in125 sp62 3183.098862
Rwpos125_63 in125 sp63 11140.846016
Rwpos125_64 in125 sp64 3183.098862
Rwpos125_65 in125 sp65 3183.098862
Rwpos125_66 in125 sp66 11140.846016
Rwpos125_67 in125 sp67 11140.846016
Rwpos125_68 in125 sp68 11140.846016
Rwpos125_69 in125 sp69 11140.846016
Rwpos125_70 in125 sp70 3183.098862
Rwpos125_71 in125 sp71 3183.098862
Rwpos125_72 in125 sp72 11140.846016
Rwpos125_73 in125 sp73 11140.846016
Rwpos125_74 in125 sp74 3183.098862
Rwpos125_75 in125 sp75 11140.846016
Rwpos125_76 in125 sp76 3183.098862
Rwpos125_77 in125 sp77 3183.098862
Rwpos125_78 in125 sp78 11140.846016
Rwpos125_79 in125 sp79 11140.846016
Rwpos125_80 in125 sp80 11140.846016
Rwpos125_81 in125 sp81 3183.098862
Rwpos125_82 in125 sp82 11140.846016
Rwpos125_83 in125 sp83 11140.846016
Rwpos125_84 in125 sp84 3183.098862
Rwpos125_85 in125 sp85 3183.098862
Rwpos125_86 in125 sp86 3183.098862
Rwpos125_87 in125 sp87 11140.846016
Rwpos125_88 in125 sp88 3183.098862
Rwpos125_89 in125 sp89 11140.846016
Rwpos125_90 in125 sp90 3183.098862
Rwpos125_91 in125 sp91 3183.098862
Rwpos125_92 in125 sp92 11140.846016
Rwpos125_93 in125 sp93 11140.846016
Rwpos125_94 in125 sp94 11140.846016
Rwpos125_95 in125 sp95 3183.098862
Rwpos125_96 in125 sp96 3183.098862
Rwpos125_97 in125 sp97 3183.098862
Rwpos125_98 in125 sp98 3183.098862
Rwpos125_99 in125 sp99 3183.098862
Rwpos125_100 in125 sp100 3183.098862
Rwpos126_1 in126 sp1 3183.098862
Rwpos126_2 in126 sp2 3183.098862
Rwpos126_3 in126 sp3 3183.098862
Rwpos126_4 in126 sp4 11140.846016
Rwpos126_5 in126 sp5 3183.098862
Rwpos126_6 in126 sp6 3183.098862
Rwpos126_7 in126 sp7 3183.098862
Rwpos126_8 in126 sp8 11140.846016
Rwpos126_9 in126 sp9 3183.098862
Rwpos126_10 in126 sp10 3183.098862
Rwpos126_11 in126 sp11 11140.846016
Rwpos126_12 in126 sp12 3183.098862
Rwpos126_13 in126 sp13 11140.846016
Rwpos126_14 in126 sp14 11140.846016
Rwpos126_15 in126 sp15 11140.846016
Rwpos126_16 in126 sp16 3183.098862
Rwpos126_17 in126 sp17 3183.098862
Rwpos126_18 in126 sp18 3183.098862
Rwpos126_19 in126 sp19 3183.098862
Rwpos126_20 in126 sp20 3183.098862
Rwpos126_21 in126 sp21 3183.098862
Rwpos126_22 in126 sp22 11140.846016
Rwpos126_23 in126 sp23 3183.098862
Rwpos126_24 in126 sp24 11140.846016
Rwpos126_25 in126 sp25 3183.098862
Rwpos126_26 in126 sp26 11140.846016
Rwpos126_27 in126 sp27 11140.846016
Rwpos126_28 in126 sp28 11140.846016
Rwpos126_29 in126 sp29 3183.098862
Rwpos126_30 in126 sp30 11140.846016
Rwpos126_31 in126 sp31 3183.098862
Rwpos126_32 in126 sp32 3183.098862
Rwpos126_33 in126 sp33 11140.846016
Rwpos126_34 in126 sp34 11140.846016
Rwpos126_35 in126 sp35 11140.846016
Rwpos126_36 in126 sp36 3183.098862
Rwpos126_37 in126 sp37 11140.846016
Rwpos126_38 in126 sp38 3183.098862
Rwpos126_39 in126 sp39 11140.846016
Rwpos126_40 in126 sp40 3183.098862
Rwpos126_41 in126 sp41 11140.846016
Rwpos126_42 in126 sp42 3183.098862
Rwpos126_43 in126 sp43 11140.846016
Rwpos126_44 in126 sp44 3183.098862


**********Negative Weighted Array****************

Rwneg1_1 in1 sn1 3183.098862
Rwneg1_2 in1 sn2 11140.846016
Rwneg1_3 in1 sn3 11140.846016
Rwneg1_4 in1 sn4 11140.846016
Rwneg1_5 in1 sn5 3183.098862
Rwneg1_6 in1 sn6 11140.846016
Rwneg1_7 in1 sn7 11140.846016
Rwneg1_8 in1 sn8 3183.098862
Rwneg1_9 in1 sn9 3183.098862
Rwneg1_10 in1 sn10 11140.846016
Rwneg1_11 in1 sn11 3183.098862
Rwneg1_12 in1 sn12 11140.846016
Rwneg1_13 in1 sn13 11140.846016
Rwneg1_14 in1 sn14 11140.846016
Rwneg1_15 in1 sn15 3183.098862
Rwneg1_16 in1 sn16 11140.846016
Rwneg1_17 in1 sn17 3183.098862
Rwneg1_18 in1 sn18 3183.098862
Rwneg1_19 in1 sn19 11140.846016
Rwneg1_20 in1 sn20 11140.846016
Rwneg1_21 in1 sn21 11140.846016
Rwneg1_22 in1 sn22 11140.846016
Rwneg1_23 in1 sn23 11140.846016
Rwneg1_24 in1 sn24 11140.846016
Rwneg1_25 in1 sn25 3183.098862
Rwneg1_26 in1 sn26 11140.846016
Rwneg1_27 in1 sn27 11140.846016
Rwneg1_28 in1 sn28 3183.098862
Rwneg1_29 in1 sn29 3183.098862
Rwneg1_30 in1 sn30 11140.846016
Rwneg1_31 in1 sn31 3183.098862
Rwneg1_32 in1 sn32 11140.846016
Rwneg1_33 in1 sn33 3183.098862
Rwneg1_34 in1 sn34 11140.846016
Rwneg1_35 in1 sn35 11140.846016
Rwneg1_36 in1 sn36 3183.098862
Rwneg1_37 in1 sn37 11140.846016
Rwneg1_38 in1 sn38 11140.846016
Rwneg1_39 in1 sn39 3183.098862
Rwneg1_40 in1 sn40 3183.098862
Rwneg1_41 in1 sn41 11140.846016
Rwneg1_42 in1 sn42 11140.846016
Rwneg1_43 in1 sn43 11140.846016
Rwneg1_44 in1 sn44 3183.098862
Rwneg1_45 in1 sn45 3183.098862
Rwneg1_46 in1 sn46 11140.846016
Rwneg1_47 in1 sn47 3183.098862
Rwneg1_48 in1 sn48 3183.098862
Rwneg1_49 in1 sn49 11140.846016
Rwneg1_50 in1 sn50 11140.846016
Rwneg1_51 in1 sn51 11140.846016
Rwneg1_52 in1 sn52 3183.098862
Rwneg1_53 in1 sn53 3183.098862
Rwneg1_54 in1 sn54 3183.098862
Rwneg1_55 in1 sn55 11140.846016
Rwneg1_56 in1 sn56 11140.846016
Rwneg1_57 in1 sn57 3183.098862
Rwneg1_58 in1 sn58 11140.846016
Rwneg1_59 in1 sn59 3183.098862
Rwneg1_60 in1 sn60 11140.846016
Rwneg1_61 in1 sn61 11140.846016
Rwneg1_62 in1 sn62 3183.098862
Rwneg1_63 in1 sn63 11140.846016
Rwneg1_64 in1 sn64 11140.846016
Rwneg1_65 in1 sn65 3183.098862
Rwneg1_66 in1 sn66 3183.098862
Rwneg1_67 in1 sn67 11140.846016
Rwneg1_68 in1 sn68 3183.098862
Rwneg1_69 in1 sn69 3183.098862
Rwneg1_70 in1 sn70 11140.846016
Rwneg1_71 in1 sn71 3183.098862
Rwneg1_72 in1 sn72 3183.098862
Rwneg1_73 in1 sn73 3183.098862
Rwneg1_74 in1 sn74 11140.846016
Rwneg1_75 in1 sn75 11140.846016
Rwneg1_76 in1 sn76 11140.846016
Rwneg1_77 in1 sn77 11140.846016
Rwneg1_78 in1 sn78 3183.098862
Rwneg1_79 in1 sn79 3183.098862
Rwneg1_80 in1 sn80 3183.098862
Rwneg1_81 in1 sn81 3183.098862
Rwneg1_82 in1 sn82 11140.846016
Rwneg1_83 in1 sn83 3183.098862
Rwneg1_84 in1 sn84 3183.098862
Rwneg1_85 in1 sn85 3183.098862
Rwneg1_86 in1 sn86 3183.098862
Rwneg1_87 in1 sn87 3183.098862
Rwneg1_88 in1 sn88 3183.098862
Rwneg1_89 in1 sn89 3183.098862
Rwneg1_90 in1 sn90 3183.098862
Rwneg1_91 in1 sn91 3183.098862
Rwneg1_92 in1 sn92 11140.846016
Rwneg1_93 in1 sn93 11140.846016
Rwneg1_94 in1 sn94 3183.098862
Rwneg1_95 in1 sn95 11140.846016
Rwneg1_96 in1 sn96 3183.098862
Rwneg1_97 in1 sn97 3183.098862
Rwneg1_98 in1 sn98 3183.098862
Rwneg1_99 in1 sn99 11140.846016
Rwneg1_100 in1 sn100 11140.846016
Rwneg2_1 in2 sn1 11140.846016
Rwneg2_2 in2 sn2 11140.846016
Rwneg2_3 in2 sn3 3183.098862
Rwneg2_4 in2 sn4 11140.846016
Rwneg2_5 in2 sn5 11140.846016
Rwneg2_6 in2 sn6 3183.098862
Rwneg2_7 in2 sn7 3183.098862
Rwneg2_8 in2 sn8 11140.846016
Rwneg2_9 in2 sn9 3183.098862
Rwneg2_10 in2 sn10 11140.846016
Rwneg2_11 in2 sn11 11140.846016
Rwneg2_12 in2 sn12 11140.846016
Rwneg2_13 in2 sn13 3183.098862
Rwneg2_14 in2 sn14 11140.846016
Rwneg2_15 in2 sn15 3183.098862
Rwneg2_16 in2 sn16 3183.098862
Rwneg2_17 in2 sn17 11140.846016
Rwneg2_18 in2 sn18 11140.846016
Rwneg2_19 in2 sn19 3183.098862
Rwneg2_20 in2 sn20 3183.098862
Rwneg2_21 in2 sn21 11140.846016
Rwneg2_22 in2 sn22 11140.846016
Rwneg2_23 in2 sn23 3183.098862
Rwneg2_24 in2 sn24 3183.098862
Rwneg2_25 in2 sn25 11140.846016
Rwneg2_26 in2 sn26 3183.098862
Rwneg2_27 in2 sn27 11140.846016
Rwneg2_28 in2 sn28 11140.846016
Rwneg2_29 in2 sn29 3183.098862
Rwneg2_30 in2 sn30 11140.846016
Rwneg2_31 in2 sn31 11140.846016
Rwneg2_32 in2 sn32 11140.846016
Rwneg2_33 in2 sn33 11140.846016
Rwneg2_34 in2 sn34 11140.846016
Rwneg2_35 in2 sn35 11140.846016
Rwneg2_36 in2 sn36 3183.098862
Rwneg2_37 in2 sn37 3183.098862
Rwneg2_38 in2 sn38 3183.098862
Rwneg2_39 in2 sn39 11140.846016
Rwneg2_40 in2 sn40 11140.846016
Rwneg2_41 in2 sn41 3183.098862
Rwneg2_42 in2 sn42 3183.098862
Rwneg2_43 in2 sn43 11140.846016
Rwneg2_44 in2 sn44 3183.098862
Rwneg2_45 in2 sn45 3183.098862
Rwneg2_46 in2 sn46 11140.846016
Rwneg2_47 in2 sn47 3183.098862
Rwneg2_48 in2 sn48 3183.098862
Rwneg2_49 in2 sn49 11140.846016
Rwneg2_50 in2 sn50 3183.098862
Rwneg2_51 in2 sn51 11140.846016
Rwneg2_52 in2 sn52 3183.098862
Rwneg2_53 in2 sn53 3183.098862
Rwneg2_54 in2 sn54 11140.846016
Rwneg2_55 in2 sn55 11140.846016
Rwneg2_56 in2 sn56 3183.098862
Rwneg2_57 in2 sn57 3183.098862
Rwneg2_58 in2 sn58 11140.846016
Rwneg2_59 in2 sn59 3183.098862
Rwneg2_60 in2 sn60 3183.098862
Rwneg2_61 in2 sn61 3183.098862
Rwneg2_62 in2 sn62 3183.098862
Rwneg2_63 in2 sn63 3183.098862
Rwneg2_64 in2 sn64 3183.098862
Rwneg2_65 in2 sn65 11140.846016
Rwneg2_66 in2 sn66 3183.098862
Rwneg2_67 in2 sn67 3183.098862
Rwneg2_68 in2 sn68 3183.098862
Rwneg2_69 in2 sn69 3183.098862
Rwneg2_70 in2 sn70 3183.098862
Rwneg2_71 in2 sn71 11140.846016
Rwneg2_72 in2 sn72 3183.098862
Rwneg2_73 in2 sn73 3183.098862
Rwneg2_74 in2 sn74 3183.098862
Rwneg2_75 in2 sn75 3183.098862
Rwneg2_76 in2 sn76 3183.098862
Rwneg2_77 in2 sn77 11140.846016
Rwneg2_78 in2 sn78 11140.846016
Rwneg2_79 in2 sn79 3183.098862
Rwneg2_80 in2 sn80 11140.846016
Rwneg2_81 in2 sn81 11140.846016
Rwneg2_82 in2 sn82 3183.098862
Rwneg2_83 in2 sn83 3183.098862
Rwneg2_84 in2 sn84 11140.846016
Rwneg2_85 in2 sn85 11140.846016
Rwneg2_86 in2 sn86 3183.098862
Rwneg2_87 in2 sn87 3183.098862
Rwneg2_88 in2 sn88 3183.098862
Rwneg2_89 in2 sn89 11140.846016
Rwneg2_90 in2 sn90 3183.098862
Rwneg2_91 in2 sn91 11140.846016
Rwneg2_92 in2 sn92 11140.846016
Rwneg2_93 in2 sn93 11140.846016
Rwneg2_94 in2 sn94 11140.846016
Rwneg2_95 in2 sn95 3183.098862
Rwneg2_96 in2 sn96 11140.846016
Rwneg2_97 in2 sn97 3183.098862
Rwneg2_98 in2 sn98 3183.098862
Rwneg2_99 in2 sn99 3183.098862
Rwneg2_100 in2 sn100 3183.098862
Rwneg3_1 in3 sn1 11140.846016
Rwneg3_2 in3 sn2 3183.098862
Rwneg3_3 in3 sn3 3183.098862
Rwneg3_4 in3 sn4 11140.846016
Rwneg3_5 in3 sn5 3183.098862
Rwneg3_6 in3 sn6 3183.098862
Rwneg3_7 in3 sn7 11140.846016
Rwneg3_8 in3 sn8 3183.098862
Rwneg3_9 in3 sn9 3183.098862
Rwneg3_10 in3 sn10 3183.098862
Rwneg3_11 in3 sn11 3183.098862
Rwneg3_12 in3 sn12 11140.846016
Rwneg3_13 in3 sn13 11140.846016
Rwneg3_14 in3 sn14 3183.098862
Rwneg3_15 in3 sn15 11140.846016
Rwneg3_16 in3 sn16 11140.846016
Rwneg3_17 in3 sn17 11140.846016
Rwneg3_18 in3 sn18 11140.846016
Rwneg3_19 in3 sn19 11140.846016
Rwneg3_20 in3 sn20 3183.098862
Rwneg3_21 in3 sn21 11140.846016
Rwneg3_22 in3 sn22 11140.846016
Rwneg3_23 in3 sn23 11140.846016
Rwneg3_24 in3 sn24 3183.098862
Rwneg3_25 in3 sn25 3183.098862
Rwneg3_26 in3 sn26 3183.098862
Rwneg3_27 in3 sn27 3183.098862
Rwneg3_28 in3 sn28 3183.098862
Rwneg3_29 in3 sn29 3183.098862
Rwneg3_30 in3 sn30 11140.846016
Rwneg3_31 in3 sn31 3183.098862
Rwneg3_32 in3 sn32 11140.846016
Rwneg3_33 in3 sn33 11140.846016
Rwneg3_34 in3 sn34 11140.846016
Rwneg3_35 in3 sn35 3183.098862
Rwneg3_36 in3 sn36 11140.846016
Rwneg3_37 in3 sn37 3183.098862
Rwneg3_38 in3 sn38 3183.098862
Rwneg3_39 in3 sn39 3183.098862
Rwneg3_40 in3 sn40 11140.846016
Rwneg3_41 in3 sn41 3183.098862
Rwneg3_42 in3 sn42 3183.098862
Rwneg3_43 in3 sn43 11140.846016
Rwneg3_44 in3 sn44 3183.098862
Rwneg3_45 in3 sn45 11140.846016
Rwneg3_46 in3 sn46 3183.098862
Rwneg3_47 in3 sn47 11140.846016
Rwneg3_48 in3 sn48 3183.098862
Rwneg3_49 in3 sn49 11140.846016
Rwneg3_50 in3 sn50 3183.098862
Rwneg3_51 in3 sn51 11140.846016
Rwneg3_52 in3 sn52 3183.098862
Rwneg3_53 in3 sn53 11140.846016
Rwneg3_54 in3 sn54 11140.846016
Rwneg3_55 in3 sn55 3183.098862
Rwneg3_56 in3 sn56 3183.098862
Rwneg3_57 in3 sn57 11140.846016
Rwneg3_58 in3 sn58 3183.098862
Rwneg3_59 in3 sn59 11140.846016
Rwneg3_60 in3 sn60 3183.098862
Rwneg3_61 in3 sn61 11140.846016
Rwneg3_62 in3 sn62 3183.098862
Rwneg3_63 in3 sn63 11140.846016
Rwneg3_64 in3 sn64 3183.098862
Rwneg3_65 in3 sn65 11140.846016
Rwneg3_66 in3 sn66 11140.846016
Rwneg3_67 in3 sn67 11140.846016
Rwneg3_68 in3 sn68 3183.098862
Rwneg3_69 in3 sn69 11140.846016
Rwneg3_70 in3 sn70 11140.846016
Rwneg3_71 in3 sn71 11140.846016
Rwneg3_72 in3 sn72 3183.098862
Rwneg3_73 in3 sn73 11140.846016
Rwneg3_74 in3 sn74 3183.098862
Rwneg3_75 in3 sn75 11140.846016
Rwneg3_76 in3 sn76 3183.098862
Rwneg3_77 in3 sn77 3183.098862
Rwneg3_78 in3 sn78 11140.846016
Rwneg3_79 in3 sn79 3183.098862
Rwneg3_80 in3 sn80 3183.098862
Rwneg3_81 in3 sn81 3183.098862
Rwneg3_82 in3 sn82 11140.846016
Rwneg3_83 in3 sn83 11140.846016
Rwneg3_84 in3 sn84 3183.098862
Rwneg3_85 in3 sn85 11140.846016
Rwneg3_86 in3 sn86 11140.846016
Rwneg3_87 in3 sn87 3183.098862
Rwneg3_88 in3 sn88 11140.846016
Rwneg3_89 in3 sn89 3183.098862
Rwneg3_90 in3 sn90 11140.846016
Rwneg3_91 in3 sn91 11140.846016
Rwneg3_92 in3 sn92 11140.846016
Rwneg3_93 in3 sn93 3183.098862
Rwneg3_94 in3 sn94 3183.098862
Rwneg3_95 in3 sn95 11140.846016
Rwneg3_96 in3 sn96 3183.098862
Rwneg3_97 in3 sn97 3183.098862
Rwneg3_98 in3 sn98 11140.846016
Rwneg3_99 in3 sn99 11140.846016
Rwneg3_100 in3 sn100 3183.098862
Rwneg4_1 in4 sn1 11140.846016
Rwneg4_2 in4 sn2 11140.846016
Rwneg4_3 in4 sn3 3183.098862
Rwneg4_4 in4 sn4 11140.846016
Rwneg4_5 in4 sn5 11140.846016
Rwneg4_6 in4 sn6 3183.098862
Rwneg4_7 in4 sn7 3183.098862
Rwneg4_8 in4 sn8 11140.846016
Rwneg4_9 in4 sn9 3183.098862
Rwneg4_10 in4 sn10 3183.098862
Rwneg4_11 in4 sn11 11140.846016
Rwneg4_12 in4 sn12 3183.098862
Rwneg4_13 in4 sn13 3183.098862
Rwneg4_14 in4 sn14 3183.098862
Rwneg4_15 in4 sn15 11140.846016
Rwneg4_16 in4 sn16 3183.098862
Rwneg4_17 in4 sn17 11140.846016
Rwneg4_18 in4 sn18 3183.098862
Rwneg4_19 in4 sn19 11140.846016
Rwneg4_20 in4 sn20 3183.098862
Rwneg4_21 in4 sn21 3183.098862
Rwneg4_22 in4 sn22 3183.098862
Rwneg4_23 in4 sn23 3183.098862
Rwneg4_24 in4 sn24 11140.846016
Rwneg4_25 in4 sn25 3183.098862
Rwneg4_26 in4 sn26 11140.846016
Rwneg4_27 in4 sn27 11140.846016
Rwneg4_28 in4 sn28 11140.846016
Rwneg4_29 in4 sn29 3183.098862
Rwneg4_30 in4 sn30 3183.098862
Rwneg4_31 in4 sn31 11140.846016
Rwneg4_32 in4 sn32 3183.098862
Rwneg4_33 in4 sn33 11140.846016
Rwneg4_34 in4 sn34 11140.846016
Rwneg4_35 in4 sn35 3183.098862
Rwneg4_36 in4 sn36 11140.846016
Rwneg4_37 in4 sn37 11140.846016
Rwneg4_38 in4 sn38 11140.846016
Rwneg4_39 in4 sn39 11140.846016
Rwneg4_40 in4 sn40 3183.098862
Rwneg4_41 in4 sn41 3183.098862
Rwneg4_42 in4 sn42 3183.098862
Rwneg4_43 in4 sn43 11140.846016
Rwneg4_44 in4 sn44 3183.098862
Rwneg4_45 in4 sn45 3183.098862
Rwneg4_46 in4 sn46 3183.098862
Rwneg4_47 in4 sn47 11140.846016
Rwneg4_48 in4 sn48 3183.098862
Rwneg4_49 in4 sn49 11140.846016
Rwneg4_50 in4 sn50 11140.846016
Rwneg4_51 in4 sn51 11140.846016
Rwneg4_52 in4 sn52 11140.846016
Rwneg4_53 in4 sn53 11140.846016
Rwneg4_54 in4 sn54 11140.846016
Rwneg4_55 in4 sn55 3183.098862
Rwneg4_56 in4 sn56 3183.098862
Rwneg4_57 in4 sn57 3183.098862
Rwneg4_58 in4 sn58 11140.846016
Rwneg4_59 in4 sn59 3183.098862
Rwneg4_60 in4 sn60 3183.098862
Rwneg4_61 in4 sn61 11140.846016
Rwneg4_62 in4 sn62 3183.098862
Rwneg4_63 in4 sn63 3183.098862
Rwneg4_64 in4 sn64 11140.846016
Rwneg4_65 in4 sn65 11140.846016
Rwneg4_66 in4 sn66 3183.098862
Rwneg4_67 in4 sn67 3183.098862
Rwneg4_68 in4 sn68 11140.846016
Rwneg4_69 in4 sn69 11140.846016
Rwneg4_70 in4 sn70 11140.846016
Rwneg4_71 in4 sn71 3183.098862
Rwneg4_72 in4 sn72 11140.846016
Rwneg4_73 in4 sn73 11140.846016
Rwneg4_74 in4 sn74 3183.098862
Rwneg4_75 in4 sn75 3183.098862
Rwneg4_76 in4 sn76 11140.846016
Rwneg4_77 in4 sn77 3183.098862
Rwneg4_78 in4 sn78 11140.846016
Rwneg4_79 in4 sn79 3183.098862
Rwneg4_80 in4 sn80 11140.846016
Rwneg4_81 in4 sn81 11140.846016
Rwneg4_82 in4 sn82 11140.846016
Rwneg4_83 in4 sn83 3183.098862
Rwneg4_84 in4 sn84 3183.098862
Rwneg4_85 in4 sn85 3183.098862
Rwneg4_86 in4 sn86 3183.098862
Rwneg4_87 in4 sn87 11140.846016
Rwneg4_88 in4 sn88 11140.846016
Rwneg4_89 in4 sn89 11140.846016
Rwneg4_90 in4 sn90 11140.846016
Rwneg4_91 in4 sn91 11140.846016
Rwneg4_92 in4 sn92 11140.846016
Rwneg4_93 in4 sn93 3183.098862
Rwneg4_94 in4 sn94 11140.846016
Rwneg4_95 in4 sn95 11140.846016
Rwneg4_96 in4 sn96 11140.846016
Rwneg4_97 in4 sn97 3183.098862
Rwneg4_98 in4 sn98 3183.098862
Rwneg4_99 in4 sn99 11140.846016
Rwneg4_100 in4 sn100 3183.098862
Rwneg5_1 in5 sn1 3183.098862
Rwneg5_2 in5 sn2 3183.098862
Rwneg5_3 in5 sn3 11140.846016
Rwneg5_4 in5 sn4 3183.098862
Rwneg5_5 in5 sn5 11140.846016
Rwneg5_6 in5 sn6 11140.846016
Rwneg5_7 in5 sn7 3183.098862
Rwneg5_8 in5 sn8 3183.098862
Rwneg5_9 in5 sn9 11140.846016
Rwneg5_10 in5 sn10 3183.098862
Rwneg5_11 in5 sn11 3183.098862
Rwneg5_12 in5 sn12 11140.846016
Rwneg5_13 in5 sn13 11140.846016
Rwneg5_14 in5 sn14 11140.846016
Rwneg5_15 in5 sn15 3183.098862
Rwneg5_16 in5 sn16 3183.098862
Rwneg5_17 in5 sn17 11140.846016
Rwneg5_18 in5 sn18 11140.846016
Rwneg5_19 in5 sn19 3183.098862
Rwneg5_20 in5 sn20 11140.846016
Rwneg5_21 in5 sn21 11140.846016
Rwneg5_22 in5 sn22 11140.846016
Rwneg5_23 in5 sn23 11140.846016
Rwneg5_24 in5 sn24 3183.098862
Rwneg5_25 in5 sn25 11140.846016
Rwneg5_26 in5 sn26 3183.098862
Rwneg5_27 in5 sn27 11140.846016
Rwneg5_28 in5 sn28 11140.846016
Rwneg5_29 in5 sn29 3183.098862
Rwneg5_30 in5 sn30 3183.098862
Rwneg5_31 in5 sn31 3183.098862
Rwneg5_32 in5 sn32 3183.098862
Rwneg5_33 in5 sn33 3183.098862
Rwneg5_34 in5 sn34 11140.846016
Rwneg5_35 in5 sn35 3183.098862
Rwneg5_36 in5 sn36 11140.846016
Rwneg5_37 in5 sn37 3183.098862
Rwneg5_38 in5 sn38 3183.098862
Rwneg5_39 in5 sn39 11140.846016
Rwneg5_40 in5 sn40 3183.098862
Rwneg5_41 in5 sn41 3183.098862
Rwneg5_42 in5 sn42 11140.846016
Rwneg5_43 in5 sn43 3183.098862
Rwneg5_44 in5 sn44 3183.098862
Rwneg5_45 in5 sn45 11140.846016
Rwneg5_46 in5 sn46 11140.846016
Rwneg5_47 in5 sn47 11140.846016
Rwneg5_48 in5 sn48 3183.098862
Rwneg5_49 in5 sn49 11140.846016
Rwneg5_50 in5 sn50 11140.846016
Rwneg5_51 in5 sn51 3183.098862
Rwneg5_52 in5 sn52 11140.846016
Rwneg5_53 in5 sn53 11140.846016
Rwneg5_54 in5 sn54 3183.098862
Rwneg5_55 in5 sn55 11140.846016
Rwneg5_56 in5 sn56 11140.846016
Rwneg5_57 in5 sn57 11140.846016
Rwneg5_58 in5 sn58 11140.846016
Rwneg5_59 in5 sn59 3183.098862
Rwneg5_60 in5 sn60 11140.846016
Rwneg5_61 in5 sn61 3183.098862
Rwneg5_62 in5 sn62 11140.846016
Rwneg5_63 in5 sn63 3183.098862
Rwneg5_64 in5 sn64 3183.098862
Rwneg5_65 in5 sn65 3183.098862
Rwneg5_66 in5 sn66 11140.846016
Rwneg5_67 in5 sn67 11140.846016
Rwneg5_68 in5 sn68 11140.846016
Rwneg5_69 in5 sn69 11140.846016
Rwneg5_70 in5 sn70 11140.846016
Rwneg5_71 in5 sn71 3183.098862
Rwneg5_72 in5 sn72 3183.098862
Rwneg5_73 in5 sn73 11140.846016
Rwneg5_74 in5 sn74 11140.846016
Rwneg5_75 in5 sn75 11140.846016
Rwneg5_76 in5 sn76 3183.098862
Rwneg5_77 in5 sn77 11140.846016
Rwneg5_78 in5 sn78 11140.846016
Rwneg5_79 in5 sn79 3183.098862
Rwneg5_80 in5 sn80 11140.846016
Rwneg5_81 in5 sn81 3183.098862
Rwneg5_82 in5 sn82 3183.098862
Rwneg5_83 in5 sn83 11140.846016
Rwneg5_84 in5 sn84 3183.098862
Rwneg5_85 in5 sn85 11140.846016
Rwneg5_86 in5 sn86 11140.846016
Rwneg5_87 in5 sn87 3183.098862
Rwneg5_88 in5 sn88 3183.098862
Rwneg5_89 in5 sn89 11140.846016
Rwneg5_90 in5 sn90 3183.098862
Rwneg5_91 in5 sn91 11140.846016
Rwneg5_92 in5 sn92 11140.846016
Rwneg5_93 in5 sn93 11140.846016
Rwneg5_94 in5 sn94 3183.098862
Rwneg5_95 in5 sn95 11140.846016
Rwneg5_96 in5 sn96 3183.098862
Rwneg5_97 in5 sn97 11140.846016
Rwneg5_98 in5 sn98 3183.098862
Rwneg5_99 in5 sn99 3183.098862
Rwneg5_100 in5 sn100 11140.846016
Rwneg6_1 in6 sn1 3183.098862
Rwneg6_2 in6 sn2 3183.098862
Rwneg6_3 in6 sn3 11140.846016
Rwneg6_4 in6 sn4 11140.846016
Rwneg6_5 in6 sn5 11140.846016
Rwneg6_6 in6 sn6 3183.098862
Rwneg6_7 in6 sn7 11140.846016
Rwneg6_8 in6 sn8 3183.098862
Rwneg6_9 in6 sn9 3183.098862
Rwneg6_10 in6 sn10 3183.098862
Rwneg6_11 in6 sn11 11140.846016
Rwneg6_12 in6 sn12 3183.098862
Rwneg6_13 in6 sn13 11140.846016
Rwneg6_14 in6 sn14 11140.846016
Rwneg6_15 in6 sn15 3183.098862
Rwneg6_16 in6 sn16 11140.846016
Rwneg6_17 in6 sn17 11140.846016
Rwneg6_18 in6 sn18 11140.846016
Rwneg6_19 in6 sn19 11140.846016
Rwneg6_20 in6 sn20 11140.846016
Rwneg6_21 in6 sn21 11140.846016
Rwneg6_22 in6 sn22 3183.098862
Rwneg6_23 in6 sn23 3183.098862
Rwneg6_24 in6 sn24 3183.098862
Rwneg6_25 in6 sn25 11140.846016
Rwneg6_26 in6 sn26 3183.098862
Rwneg6_27 in6 sn27 11140.846016
Rwneg6_28 in6 sn28 3183.098862
Rwneg6_29 in6 sn29 11140.846016
Rwneg6_30 in6 sn30 11140.846016
Rwneg6_31 in6 sn31 11140.846016
Rwneg6_32 in6 sn32 3183.098862
Rwneg6_33 in6 sn33 11140.846016
Rwneg6_34 in6 sn34 3183.098862
Rwneg6_35 in6 sn35 11140.846016
Rwneg6_36 in6 sn36 11140.846016
Rwneg6_37 in6 sn37 11140.846016
Rwneg6_38 in6 sn38 11140.846016
Rwneg6_39 in6 sn39 11140.846016
Rwneg6_40 in6 sn40 11140.846016
Rwneg6_41 in6 sn41 3183.098862
Rwneg6_42 in6 sn42 11140.846016
Rwneg6_43 in6 sn43 11140.846016
Rwneg6_44 in6 sn44 3183.098862
Rwneg6_45 in6 sn45 3183.098862
Rwneg6_46 in6 sn46 3183.098862
Rwneg6_47 in6 sn47 3183.098862
Rwneg6_48 in6 sn48 11140.846016
Rwneg6_49 in6 sn49 3183.098862
Rwneg6_50 in6 sn50 3183.098862
Rwneg6_51 in6 sn51 11140.846016
Rwneg6_52 in6 sn52 11140.846016
Rwneg6_53 in6 sn53 11140.846016
Rwneg6_54 in6 sn54 11140.846016
Rwneg6_55 in6 sn55 11140.846016
Rwneg6_56 in6 sn56 11140.846016
Rwneg6_57 in6 sn57 3183.098862
Rwneg6_58 in6 sn58 11140.846016
Rwneg6_59 in6 sn59 3183.098862
Rwneg6_60 in6 sn60 3183.098862
Rwneg6_61 in6 sn61 11140.846016
Rwneg6_62 in6 sn62 11140.846016
Rwneg6_63 in6 sn63 11140.846016
Rwneg6_64 in6 sn64 3183.098862
Rwneg6_65 in6 sn65 11140.846016
Rwneg6_66 in6 sn66 11140.846016
Rwneg6_67 in6 sn67 11140.846016
Rwneg6_68 in6 sn68 3183.098862
Rwneg6_69 in6 sn69 3183.098862
Rwneg6_70 in6 sn70 11140.846016
Rwneg6_71 in6 sn71 3183.098862
Rwneg6_72 in6 sn72 11140.846016
Rwneg6_73 in6 sn73 11140.846016
Rwneg6_74 in6 sn74 3183.098862
Rwneg6_75 in6 sn75 11140.846016
Rwneg6_76 in6 sn76 3183.098862
Rwneg6_77 in6 sn77 3183.098862
Rwneg6_78 in6 sn78 11140.846016
Rwneg6_79 in6 sn79 11140.846016
Rwneg6_80 in6 sn80 11140.846016
Rwneg6_81 in6 sn81 11140.846016
Rwneg6_82 in6 sn82 3183.098862
Rwneg6_83 in6 sn83 11140.846016
Rwneg6_84 in6 sn84 11140.846016
Rwneg6_85 in6 sn85 3183.098862
Rwneg6_86 in6 sn86 11140.846016
Rwneg6_87 in6 sn87 3183.098862
Rwneg6_88 in6 sn88 11140.846016
Rwneg6_89 in6 sn89 3183.098862
Rwneg6_90 in6 sn90 11140.846016
Rwneg6_91 in6 sn91 11140.846016
Rwneg6_92 in6 sn92 11140.846016
Rwneg6_93 in6 sn93 11140.846016
Rwneg6_94 in6 sn94 11140.846016
Rwneg6_95 in6 sn95 11140.846016
Rwneg6_96 in6 sn96 3183.098862
Rwneg6_97 in6 sn97 3183.098862
Rwneg6_98 in6 sn98 3183.098862
Rwneg6_99 in6 sn99 3183.098862
Rwneg6_100 in6 sn100 11140.846016
Rwneg7_1 in7 sn1 11140.846016
Rwneg7_2 in7 sn2 11140.846016
Rwneg7_3 in7 sn3 3183.098862
Rwneg7_4 in7 sn4 11140.846016
Rwneg7_5 in7 sn5 3183.098862
Rwneg7_6 in7 sn6 3183.098862
Rwneg7_7 in7 sn7 11140.846016
Rwneg7_8 in7 sn8 11140.846016
Rwneg7_9 in7 sn9 11140.846016
Rwneg7_10 in7 sn10 3183.098862
Rwneg7_11 in7 sn11 11140.846016
Rwneg7_12 in7 sn12 11140.846016
Rwneg7_13 in7 sn13 3183.098862
Rwneg7_14 in7 sn14 3183.098862
Rwneg7_15 in7 sn15 3183.098862
Rwneg7_16 in7 sn16 11140.846016
Rwneg7_17 in7 sn17 3183.098862
Rwneg7_18 in7 sn18 11140.846016
Rwneg7_19 in7 sn19 11140.846016
Rwneg7_20 in7 sn20 3183.098862
Rwneg7_21 in7 sn21 3183.098862
Rwneg7_22 in7 sn22 3183.098862
Rwneg7_23 in7 sn23 3183.098862
Rwneg7_24 in7 sn24 11140.846016
Rwneg7_25 in7 sn25 3183.098862
Rwneg7_26 in7 sn26 3183.098862
Rwneg7_27 in7 sn27 11140.846016
Rwneg7_28 in7 sn28 11140.846016
Rwneg7_29 in7 sn29 3183.098862
Rwneg7_30 in7 sn30 11140.846016
Rwneg7_31 in7 sn31 11140.846016
Rwneg7_32 in7 sn32 3183.098862
Rwneg7_33 in7 sn33 11140.846016
Rwneg7_34 in7 sn34 11140.846016
Rwneg7_35 in7 sn35 11140.846016
Rwneg7_36 in7 sn36 3183.098862
Rwneg7_37 in7 sn37 11140.846016
Rwneg7_38 in7 sn38 11140.846016
Rwneg7_39 in7 sn39 3183.098862
Rwneg7_40 in7 sn40 11140.846016
Rwneg7_41 in7 sn41 3183.098862
Rwneg7_42 in7 sn42 3183.098862
Rwneg7_43 in7 sn43 3183.098862
Rwneg7_44 in7 sn44 3183.098862
Rwneg7_45 in7 sn45 11140.846016
Rwneg7_46 in7 sn46 3183.098862
Rwneg7_47 in7 sn47 11140.846016
Rwneg7_48 in7 sn48 3183.098862
Rwneg7_49 in7 sn49 3183.098862
Rwneg7_50 in7 sn50 3183.098862
Rwneg7_51 in7 sn51 3183.098862
Rwneg7_52 in7 sn52 11140.846016
Rwneg7_53 in7 sn53 3183.098862
Rwneg7_54 in7 sn54 3183.098862
Rwneg7_55 in7 sn55 3183.098862
Rwneg7_56 in7 sn56 3183.098862
Rwneg7_57 in7 sn57 11140.846016
Rwneg7_58 in7 sn58 11140.846016
Rwneg7_59 in7 sn59 3183.098862
Rwneg7_60 in7 sn60 3183.098862
Rwneg7_61 in7 sn61 11140.846016
Rwneg7_62 in7 sn62 3183.098862
Rwneg7_63 in7 sn63 11140.846016
Rwneg7_64 in7 sn64 11140.846016
Rwneg7_65 in7 sn65 11140.846016
Rwneg7_66 in7 sn66 11140.846016
Rwneg7_67 in7 sn67 3183.098862
Rwneg7_68 in7 sn68 11140.846016
Rwneg7_69 in7 sn69 11140.846016
Rwneg7_70 in7 sn70 3183.098862
Rwneg7_71 in7 sn71 3183.098862
Rwneg7_72 in7 sn72 3183.098862
Rwneg7_73 in7 sn73 11140.846016
Rwneg7_74 in7 sn74 3183.098862
Rwneg7_75 in7 sn75 3183.098862
Rwneg7_76 in7 sn76 3183.098862
Rwneg7_77 in7 sn77 3183.098862
Rwneg7_78 in7 sn78 3183.098862
Rwneg7_79 in7 sn79 3183.098862
Rwneg7_80 in7 sn80 11140.846016
Rwneg7_81 in7 sn81 3183.098862
Rwneg7_82 in7 sn82 11140.846016
Rwneg7_83 in7 sn83 3183.098862
Rwneg7_84 in7 sn84 11140.846016
Rwneg7_85 in7 sn85 11140.846016
Rwneg7_86 in7 sn86 3183.098862
Rwneg7_87 in7 sn87 3183.098862
Rwneg7_88 in7 sn88 3183.098862
Rwneg7_89 in7 sn89 11140.846016
Rwneg7_90 in7 sn90 3183.098862
Rwneg7_91 in7 sn91 11140.846016
Rwneg7_92 in7 sn92 11140.846016
Rwneg7_93 in7 sn93 3183.098862
Rwneg7_94 in7 sn94 3183.098862
Rwneg7_95 in7 sn95 11140.846016
Rwneg7_96 in7 sn96 11140.846016
Rwneg7_97 in7 sn97 11140.846016
Rwneg7_98 in7 sn98 11140.846016
Rwneg7_99 in7 sn99 3183.098862
Rwneg7_100 in7 sn100 11140.846016
Rwneg8_1 in8 sn1 11140.846016
Rwneg8_2 in8 sn2 3183.098862
Rwneg8_3 in8 sn3 3183.098862
Rwneg8_4 in8 sn4 11140.846016
Rwneg8_5 in8 sn5 3183.098862
Rwneg8_6 in8 sn6 3183.098862
Rwneg8_7 in8 sn7 3183.098862
Rwneg8_8 in8 sn8 3183.098862
Rwneg8_9 in8 sn9 11140.846016
Rwneg8_10 in8 sn10 11140.846016
Rwneg8_11 in8 sn11 3183.098862
Rwneg8_12 in8 sn12 11140.846016
Rwneg8_13 in8 sn13 3183.098862
Rwneg8_14 in8 sn14 11140.846016
Rwneg8_15 in8 sn15 3183.098862
Rwneg8_16 in8 sn16 11140.846016
Rwneg8_17 in8 sn17 3183.098862
Rwneg8_18 in8 sn18 3183.098862
Rwneg8_19 in8 sn19 11140.846016
Rwneg8_20 in8 sn20 3183.098862
Rwneg8_21 in8 sn21 11140.846016
Rwneg8_22 in8 sn22 3183.098862
Rwneg8_23 in8 sn23 11140.846016
Rwneg8_24 in8 sn24 3183.098862
Rwneg8_25 in8 sn25 3183.098862
Rwneg8_26 in8 sn26 11140.846016
Rwneg8_27 in8 sn27 3183.098862
Rwneg8_28 in8 sn28 11140.846016
Rwneg8_29 in8 sn29 11140.846016
Rwneg8_30 in8 sn30 3183.098862
Rwneg8_31 in8 sn31 3183.098862
Rwneg8_32 in8 sn32 11140.846016
Rwneg8_33 in8 sn33 11140.846016
Rwneg8_34 in8 sn34 11140.846016
Rwneg8_35 in8 sn35 3183.098862
Rwneg8_36 in8 sn36 11140.846016
Rwneg8_37 in8 sn37 3183.098862
Rwneg8_38 in8 sn38 11140.846016
Rwneg8_39 in8 sn39 11140.846016
Rwneg8_40 in8 sn40 3183.098862
Rwneg8_41 in8 sn41 11140.846016
Rwneg8_42 in8 sn42 11140.846016
Rwneg8_43 in8 sn43 11140.846016
Rwneg8_44 in8 sn44 3183.098862
Rwneg8_45 in8 sn45 11140.846016
Rwneg8_46 in8 sn46 11140.846016
Rwneg8_47 in8 sn47 11140.846016
Rwneg8_48 in8 sn48 11140.846016
Rwneg8_49 in8 sn49 3183.098862
Rwneg8_50 in8 sn50 11140.846016
Rwneg8_51 in8 sn51 3183.098862
Rwneg8_52 in8 sn52 3183.098862
Rwneg8_53 in8 sn53 11140.846016
Rwneg8_54 in8 sn54 3183.098862
Rwneg8_55 in8 sn55 3183.098862
Rwneg8_56 in8 sn56 11140.846016
Rwneg8_57 in8 sn57 3183.098862
Rwneg8_58 in8 sn58 3183.098862
Rwneg8_59 in8 sn59 3183.098862
Rwneg8_60 in8 sn60 3183.098862
Rwneg8_61 in8 sn61 11140.846016
Rwneg8_62 in8 sn62 11140.846016
Rwneg8_63 in8 sn63 11140.846016
Rwneg8_64 in8 sn64 11140.846016
Rwneg8_65 in8 sn65 3183.098862
Rwneg8_66 in8 sn66 11140.846016
Rwneg8_67 in8 sn67 3183.098862
Rwneg8_68 in8 sn68 11140.846016
Rwneg8_69 in8 sn69 11140.846016
Rwneg8_70 in8 sn70 11140.846016
Rwneg8_71 in8 sn71 3183.098862
Rwneg8_72 in8 sn72 3183.098862
Rwneg8_73 in8 sn73 11140.846016
Rwneg8_74 in8 sn74 3183.098862
Rwneg8_75 in8 sn75 3183.098862
Rwneg8_76 in8 sn76 3183.098862
Rwneg8_77 in8 sn77 11140.846016
Rwneg8_78 in8 sn78 11140.846016
Rwneg8_79 in8 sn79 3183.098862
Rwneg8_80 in8 sn80 3183.098862
Rwneg8_81 in8 sn81 3183.098862
Rwneg8_82 in8 sn82 11140.846016
Rwneg8_83 in8 sn83 11140.846016
Rwneg8_84 in8 sn84 3183.098862
Rwneg8_85 in8 sn85 3183.098862
Rwneg8_86 in8 sn86 3183.098862
Rwneg8_87 in8 sn87 3183.098862
Rwneg8_88 in8 sn88 11140.846016
Rwneg8_89 in8 sn89 11140.846016
Rwneg8_90 in8 sn90 3183.098862
Rwneg8_91 in8 sn91 3183.098862
Rwneg8_92 in8 sn92 11140.846016
Rwneg8_93 in8 sn93 3183.098862
Rwneg8_94 in8 sn94 11140.846016
Rwneg8_95 in8 sn95 11140.846016
Rwneg8_96 in8 sn96 3183.098862
Rwneg8_97 in8 sn97 3183.098862
Rwneg8_98 in8 sn98 3183.098862
Rwneg8_99 in8 sn99 3183.098862
Rwneg8_100 in8 sn100 3183.098862
Rwneg9_1 in9 sn1 3183.098862
Rwneg9_2 in9 sn2 3183.098862
Rwneg9_3 in9 sn3 3183.098862
Rwneg9_4 in9 sn4 11140.846016
Rwneg9_5 in9 sn5 3183.098862
Rwneg9_6 in9 sn6 11140.846016
Rwneg9_7 in9 sn7 3183.098862
Rwneg9_8 in9 sn8 3183.098862
Rwneg9_9 in9 sn9 11140.846016
Rwneg9_10 in9 sn10 3183.098862
Rwneg9_11 in9 sn11 3183.098862
Rwneg9_12 in9 sn12 3183.098862
Rwneg9_13 in9 sn13 3183.098862
Rwneg9_14 in9 sn14 3183.098862
Rwneg9_15 in9 sn15 3183.098862
Rwneg9_16 in9 sn16 11140.846016
Rwneg9_17 in9 sn17 11140.846016
Rwneg9_18 in9 sn18 11140.846016
Rwneg9_19 in9 sn19 3183.098862
Rwneg9_20 in9 sn20 3183.098862
Rwneg9_21 in9 sn21 11140.846016
Rwneg9_22 in9 sn22 3183.098862
Rwneg9_23 in9 sn23 3183.098862
Rwneg9_24 in9 sn24 11140.846016
Rwneg9_25 in9 sn25 11140.846016
Rwneg9_26 in9 sn26 11140.846016
Rwneg9_27 in9 sn27 11140.846016
Rwneg9_28 in9 sn28 3183.098862
Rwneg9_29 in9 sn29 11140.846016
Rwneg9_30 in9 sn30 3183.098862
Rwneg9_31 in9 sn31 11140.846016
Rwneg9_32 in9 sn32 3183.098862
Rwneg9_33 in9 sn33 11140.846016
Rwneg9_34 in9 sn34 3183.098862
Rwneg9_35 in9 sn35 3183.098862
Rwneg9_36 in9 sn36 3183.098862
Rwneg9_37 in9 sn37 11140.846016
Rwneg9_38 in9 sn38 3183.098862
Rwneg9_39 in9 sn39 11140.846016
Rwneg9_40 in9 sn40 11140.846016
Rwneg9_41 in9 sn41 11140.846016
Rwneg9_42 in9 sn42 3183.098862
Rwneg9_43 in9 sn43 3183.098862
Rwneg9_44 in9 sn44 11140.846016
Rwneg9_45 in9 sn45 3183.098862
Rwneg9_46 in9 sn46 3183.098862
Rwneg9_47 in9 sn47 11140.846016
Rwneg9_48 in9 sn48 3183.098862
Rwneg9_49 in9 sn49 3183.098862
Rwneg9_50 in9 sn50 3183.098862
Rwneg9_51 in9 sn51 3183.098862
Rwneg9_52 in9 sn52 11140.846016
Rwneg9_53 in9 sn53 11140.846016
Rwneg9_54 in9 sn54 3183.098862
Rwneg9_55 in9 sn55 3183.098862
Rwneg9_56 in9 sn56 11140.846016
Rwneg9_57 in9 sn57 3183.098862
Rwneg9_58 in9 sn58 11140.846016
Rwneg9_59 in9 sn59 3183.098862
Rwneg9_60 in9 sn60 3183.098862
Rwneg9_61 in9 sn61 11140.846016
Rwneg9_62 in9 sn62 3183.098862
Rwneg9_63 in9 sn63 11140.846016
Rwneg9_64 in9 sn64 11140.846016
Rwneg9_65 in9 sn65 11140.846016
Rwneg9_66 in9 sn66 3183.098862
Rwneg9_67 in9 sn67 11140.846016
Rwneg9_68 in9 sn68 3183.098862
Rwneg9_69 in9 sn69 11140.846016
Rwneg9_70 in9 sn70 3183.098862
Rwneg9_71 in9 sn71 3183.098862
Rwneg9_72 in9 sn72 3183.098862
Rwneg9_73 in9 sn73 3183.098862
Rwneg9_74 in9 sn74 11140.846016
Rwneg9_75 in9 sn75 11140.846016
Rwneg9_76 in9 sn76 3183.098862
Rwneg9_77 in9 sn77 11140.846016
Rwneg9_78 in9 sn78 3183.098862
Rwneg9_79 in9 sn79 11140.846016
Rwneg9_80 in9 sn80 3183.098862
Rwneg9_81 in9 sn81 3183.098862
Rwneg9_82 in9 sn82 11140.846016
Rwneg9_83 in9 sn83 11140.846016
Rwneg9_84 in9 sn84 3183.098862
Rwneg9_85 in9 sn85 11140.846016
Rwneg9_86 in9 sn86 3183.098862
Rwneg9_87 in9 sn87 3183.098862
Rwneg9_88 in9 sn88 11140.846016
Rwneg9_89 in9 sn89 11140.846016
Rwneg9_90 in9 sn90 3183.098862
Rwneg9_91 in9 sn91 11140.846016
Rwneg9_92 in9 sn92 11140.846016
Rwneg9_93 in9 sn93 3183.098862
Rwneg9_94 in9 sn94 11140.846016
Rwneg9_95 in9 sn95 11140.846016
Rwneg9_96 in9 sn96 3183.098862
Rwneg9_97 in9 sn97 3183.098862
Rwneg9_98 in9 sn98 11140.846016
Rwneg9_99 in9 sn99 3183.098862
Rwneg9_100 in9 sn100 11140.846016
Rwneg10_1 in10 sn1 3183.098862
Rwneg10_2 in10 sn2 3183.098862
Rwneg10_3 in10 sn3 3183.098862
Rwneg10_4 in10 sn4 11140.846016
Rwneg10_5 in10 sn5 3183.098862
Rwneg10_6 in10 sn6 3183.098862
Rwneg10_7 in10 sn7 3183.098862
Rwneg10_8 in10 sn8 3183.098862
Rwneg10_9 in10 sn9 11140.846016
Rwneg10_10 in10 sn10 11140.846016
Rwneg10_11 in10 sn11 11140.846016
Rwneg10_12 in10 sn12 3183.098862
Rwneg10_13 in10 sn13 11140.846016
Rwneg10_14 in10 sn14 3183.098862
Rwneg10_15 in10 sn15 3183.098862
Rwneg10_16 in10 sn16 3183.098862
Rwneg10_17 in10 sn17 3183.098862
Rwneg10_18 in10 sn18 3183.098862
Rwneg10_19 in10 sn19 3183.098862
Rwneg10_20 in10 sn20 3183.098862
Rwneg10_21 in10 sn21 11140.846016
Rwneg10_22 in10 sn22 11140.846016
Rwneg10_23 in10 sn23 11140.846016
Rwneg10_24 in10 sn24 11140.846016
Rwneg10_25 in10 sn25 3183.098862
Rwneg10_26 in10 sn26 11140.846016
Rwneg10_27 in10 sn27 3183.098862
Rwneg10_28 in10 sn28 3183.098862
Rwneg10_29 in10 sn29 11140.846016
Rwneg10_30 in10 sn30 3183.098862
Rwneg10_31 in10 sn31 3183.098862
Rwneg10_32 in10 sn32 3183.098862
Rwneg10_33 in10 sn33 3183.098862
Rwneg10_34 in10 sn34 11140.846016
Rwneg10_35 in10 sn35 3183.098862
Rwneg10_36 in10 sn36 11140.846016
Rwneg10_37 in10 sn37 11140.846016
Rwneg10_38 in10 sn38 11140.846016
Rwneg10_39 in10 sn39 11140.846016
Rwneg10_40 in10 sn40 3183.098862
Rwneg10_41 in10 sn41 3183.098862
Rwneg10_42 in10 sn42 3183.098862
Rwneg10_43 in10 sn43 11140.846016
Rwneg10_44 in10 sn44 11140.846016
Rwneg10_45 in10 sn45 3183.098862
Rwneg10_46 in10 sn46 11140.846016
Rwneg10_47 in10 sn47 11140.846016
Rwneg10_48 in10 sn48 11140.846016
Rwneg10_49 in10 sn49 3183.098862
Rwneg10_50 in10 sn50 11140.846016
Rwneg10_51 in10 sn51 3183.098862
Rwneg10_52 in10 sn52 11140.846016
Rwneg10_53 in10 sn53 3183.098862
Rwneg10_54 in10 sn54 3183.098862
Rwneg10_55 in10 sn55 3183.098862
Rwneg10_56 in10 sn56 3183.098862
Rwneg10_57 in10 sn57 3183.098862
Rwneg10_58 in10 sn58 3183.098862
Rwneg10_59 in10 sn59 11140.846016
Rwneg10_60 in10 sn60 11140.846016
Rwneg10_61 in10 sn61 3183.098862
Rwneg10_62 in10 sn62 11140.846016
Rwneg10_63 in10 sn63 11140.846016
Rwneg10_64 in10 sn64 3183.098862
Rwneg10_65 in10 sn65 3183.098862
Rwneg10_66 in10 sn66 3183.098862
Rwneg10_67 in10 sn67 3183.098862
Rwneg10_68 in10 sn68 3183.098862
Rwneg10_69 in10 sn69 11140.846016
Rwneg10_70 in10 sn70 3183.098862
Rwneg10_71 in10 sn71 3183.098862
Rwneg10_72 in10 sn72 3183.098862
Rwneg10_73 in10 sn73 3183.098862
Rwneg10_74 in10 sn74 11140.846016
Rwneg10_75 in10 sn75 11140.846016
Rwneg10_76 in10 sn76 11140.846016
Rwneg10_77 in10 sn77 3183.098862
Rwneg10_78 in10 sn78 3183.098862
Rwneg10_79 in10 sn79 11140.846016
Rwneg10_80 in10 sn80 3183.098862
Rwneg10_81 in10 sn81 3183.098862
Rwneg10_82 in10 sn82 3183.098862
Rwneg10_83 in10 sn83 11140.846016
Rwneg10_84 in10 sn84 3183.098862
Rwneg10_85 in10 sn85 11140.846016
Rwneg10_86 in10 sn86 11140.846016
Rwneg10_87 in10 sn87 3183.098862
Rwneg10_88 in10 sn88 11140.846016
Rwneg10_89 in10 sn89 3183.098862
Rwneg10_90 in10 sn90 3183.098862
Rwneg10_91 in10 sn91 11140.846016
Rwneg10_92 in10 sn92 11140.846016
Rwneg10_93 in10 sn93 3183.098862
Rwneg10_94 in10 sn94 3183.098862
Rwneg10_95 in10 sn95 3183.098862
Rwneg10_96 in10 sn96 11140.846016
Rwneg10_97 in10 sn97 11140.846016
Rwneg10_98 in10 sn98 11140.846016
Rwneg10_99 in10 sn99 3183.098862
Rwneg10_100 in10 sn100 11140.846016
Rwneg11_1 in11 sn1 11140.846016
Rwneg11_2 in11 sn2 11140.846016
Rwneg11_3 in11 sn3 11140.846016
Rwneg11_4 in11 sn4 11140.846016
Rwneg11_5 in11 sn5 3183.098862
Rwneg11_6 in11 sn6 3183.098862
Rwneg11_7 in11 sn7 3183.098862
Rwneg11_8 in11 sn8 3183.098862
Rwneg11_9 in11 sn9 11140.846016
Rwneg11_10 in11 sn10 11140.846016
Rwneg11_11 in11 sn11 11140.846016
Rwneg11_12 in11 sn12 11140.846016
Rwneg11_13 in11 sn13 11140.846016
Rwneg11_14 in11 sn14 11140.846016
Rwneg11_15 in11 sn15 3183.098862
Rwneg11_16 in11 sn16 3183.098862
Rwneg11_17 in11 sn17 3183.098862
Rwneg11_18 in11 sn18 11140.846016
Rwneg11_19 in11 sn19 11140.846016
Rwneg11_20 in11 sn20 11140.846016
Rwneg11_21 in11 sn21 3183.098862
Rwneg11_22 in11 sn22 11140.846016
Rwneg11_23 in11 sn23 3183.098862
Rwneg11_24 in11 sn24 3183.098862
Rwneg11_25 in11 sn25 11140.846016
Rwneg11_26 in11 sn26 11140.846016
Rwneg11_27 in11 sn27 11140.846016
Rwneg11_28 in11 sn28 11140.846016
Rwneg11_29 in11 sn29 11140.846016
Rwneg11_30 in11 sn30 11140.846016
Rwneg11_31 in11 sn31 11140.846016
Rwneg11_32 in11 sn32 11140.846016
Rwneg11_33 in11 sn33 3183.098862
Rwneg11_34 in11 sn34 3183.098862
Rwneg11_35 in11 sn35 3183.098862
Rwneg11_36 in11 sn36 11140.846016
Rwneg11_37 in11 sn37 11140.846016
Rwneg11_38 in11 sn38 3183.098862
Rwneg11_39 in11 sn39 11140.846016
Rwneg11_40 in11 sn40 3183.098862
Rwneg11_41 in11 sn41 3183.098862
Rwneg11_42 in11 sn42 11140.846016
Rwneg11_43 in11 sn43 11140.846016
Rwneg11_44 in11 sn44 3183.098862
Rwneg11_45 in11 sn45 3183.098862
Rwneg11_46 in11 sn46 11140.846016
Rwneg11_47 in11 sn47 11140.846016
Rwneg11_48 in11 sn48 3183.098862
Rwneg11_49 in11 sn49 3183.098862
Rwneg11_50 in11 sn50 3183.098862
Rwneg11_51 in11 sn51 3183.098862
Rwneg11_52 in11 sn52 11140.846016
Rwneg11_53 in11 sn53 3183.098862
Rwneg11_54 in11 sn54 3183.098862
Rwneg11_55 in11 sn55 3183.098862
Rwneg11_56 in11 sn56 11140.846016
Rwneg11_57 in11 sn57 11140.846016
Rwneg11_58 in11 sn58 3183.098862
Rwneg11_59 in11 sn59 11140.846016
Rwneg11_60 in11 sn60 3183.098862
Rwneg11_61 in11 sn61 11140.846016
Rwneg11_62 in11 sn62 3183.098862
Rwneg11_63 in11 sn63 11140.846016
Rwneg11_64 in11 sn64 3183.098862
Rwneg11_65 in11 sn65 3183.098862
Rwneg11_66 in11 sn66 11140.846016
Rwneg11_67 in11 sn67 11140.846016
Rwneg11_68 in11 sn68 11140.846016
Rwneg11_69 in11 sn69 11140.846016
Rwneg11_70 in11 sn70 11140.846016
Rwneg11_71 in11 sn71 3183.098862
Rwneg11_72 in11 sn72 3183.098862
Rwneg11_73 in11 sn73 11140.846016
Rwneg11_74 in11 sn74 11140.846016
Rwneg11_75 in11 sn75 11140.846016
Rwneg11_76 in11 sn76 11140.846016
Rwneg11_77 in11 sn77 11140.846016
Rwneg11_78 in11 sn78 11140.846016
Rwneg11_79 in11 sn79 3183.098862
Rwneg11_80 in11 sn80 3183.098862
Rwneg11_81 in11 sn81 11140.846016
Rwneg11_82 in11 sn82 3183.098862
Rwneg11_83 in11 sn83 3183.098862
Rwneg11_84 in11 sn84 3183.098862
Rwneg11_85 in11 sn85 11140.846016
Rwneg11_86 in11 sn86 3183.098862
Rwneg11_87 in11 sn87 11140.846016
Rwneg11_88 in11 sn88 11140.846016
Rwneg11_89 in11 sn89 11140.846016
Rwneg11_90 in11 sn90 11140.846016
Rwneg11_91 in11 sn91 11140.846016
Rwneg11_92 in11 sn92 11140.846016
Rwneg11_93 in11 sn93 11140.846016
Rwneg11_94 in11 sn94 3183.098862
Rwneg11_95 in11 sn95 3183.098862
Rwneg11_96 in11 sn96 11140.846016
Rwneg11_97 in11 sn97 11140.846016
Rwneg11_98 in11 sn98 3183.098862
Rwneg11_99 in11 sn99 11140.846016
Rwneg11_100 in11 sn100 11140.846016
Rwneg12_1 in12 sn1 3183.098862
Rwneg12_2 in12 sn2 11140.846016
Rwneg12_3 in12 sn3 11140.846016
Rwneg12_4 in12 sn4 3183.098862
Rwneg12_5 in12 sn5 11140.846016
Rwneg12_6 in12 sn6 11140.846016
Rwneg12_7 in12 sn7 11140.846016
Rwneg12_8 in12 sn8 3183.098862
Rwneg12_9 in12 sn9 11140.846016
Rwneg12_10 in12 sn10 3183.098862
Rwneg12_11 in12 sn11 11140.846016
Rwneg12_12 in12 sn12 11140.846016
Rwneg12_13 in12 sn13 3183.098862
Rwneg12_14 in12 sn14 3183.098862
Rwneg12_15 in12 sn15 11140.846016
Rwneg12_16 in12 sn16 11140.846016
Rwneg12_17 in12 sn17 11140.846016
Rwneg12_18 in12 sn18 11140.846016
Rwneg12_19 in12 sn19 11140.846016
Rwneg12_20 in12 sn20 3183.098862
Rwneg12_21 in12 sn21 3183.098862
Rwneg12_22 in12 sn22 11140.846016
Rwneg12_23 in12 sn23 11140.846016
Rwneg12_24 in12 sn24 11140.846016
Rwneg12_25 in12 sn25 3183.098862
Rwneg12_26 in12 sn26 3183.098862
Rwneg12_27 in12 sn27 11140.846016
Rwneg12_28 in12 sn28 11140.846016
Rwneg12_29 in12 sn29 3183.098862
Rwneg12_30 in12 sn30 3183.098862
Rwneg12_31 in12 sn31 3183.098862
Rwneg12_32 in12 sn32 11140.846016
Rwneg12_33 in12 sn33 11140.846016
Rwneg12_34 in12 sn34 11140.846016
Rwneg12_35 in12 sn35 11140.846016
Rwneg12_36 in12 sn36 3183.098862
Rwneg12_37 in12 sn37 11140.846016
Rwneg12_38 in12 sn38 3183.098862
Rwneg12_39 in12 sn39 11140.846016
Rwneg12_40 in12 sn40 11140.846016
Rwneg12_41 in12 sn41 11140.846016
Rwneg12_42 in12 sn42 3183.098862
Rwneg12_43 in12 sn43 11140.846016
Rwneg12_44 in12 sn44 11140.846016
Rwneg12_45 in12 sn45 11140.846016
Rwneg12_46 in12 sn46 11140.846016
Rwneg12_47 in12 sn47 3183.098862
Rwneg12_48 in12 sn48 11140.846016
Rwneg12_49 in12 sn49 11140.846016
Rwneg12_50 in12 sn50 11140.846016
Rwneg12_51 in12 sn51 3183.098862
Rwneg12_52 in12 sn52 3183.098862
Rwneg12_53 in12 sn53 11140.846016
Rwneg12_54 in12 sn54 11140.846016
Rwneg12_55 in12 sn55 11140.846016
Rwneg12_56 in12 sn56 3183.098862
Rwneg12_57 in12 sn57 3183.098862
Rwneg12_58 in12 sn58 3183.098862
Rwneg12_59 in12 sn59 11140.846016
Rwneg12_60 in12 sn60 11140.846016
Rwneg12_61 in12 sn61 11140.846016
Rwneg12_62 in12 sn62 3183.098862
Rwneg12_63 in12 sn63 3183.098862
Rwneg12_64 in12 sn64 3183.098862
Rwneg12_65 in12 sn65 3183.098862
Rwneg12_66 in12 sn66 3183.098862
Rwneg12_67 in12 sn67 11140.846016
Rwneg12_68 in12 sn68 11140.846016
Rwneg12_69 in12 sn69 3183.098862
Rwneg12_70 in12 sn70 11140.846016
Rwneg12_71 in12 sn71 3183.098862
Rwneg12_72 in12 sn72 11140.846016
Rwneg12_73 in12 sn73 11140.846016
Rwneg12_74 in12 sn74 3183.098862
Rwneg12_75 in12 sn75 11140.846016
Rwneg12_76 in12 sn76 11140.846016
Rwneg12_77 in12 sn77 11140.846016
Rwneg12_78 in12 sn78 11140.846016
Rwneg12_79 in12 sn79 11140.846016
Rwneg12_80 in12 sn80 11140.846016
Rwneg12_81 in12 sn81 3183.098862
Rwneg12_82 in12 sn82 11140.846016
Rwneg12_83 in12 sn83 3183.098862
Rwneg12_84 in12 sn84 3183.098862
Rwneg12_85 in12 sn85 11140.846016
Rwneg12_86 in12 sn86 11140.846016
Rwneg12_87 in12 sn87 3183.098862
Rwneg12_88 in12 sn88 3183.098862
Rwneg12_89 in12 sn89 3183.098862
Rwneg12_90 in12 sn90 3183.098862
Rwneg12_91 in12 sn91 11140.846016
Rwneg12_92 in12 sn92 11140.846016
Rwneg12_93 in12 sn93 11140.846016
Rwneg12_94 in12 sn94 3183.098862
Rwneg12_95 in12 sn95 11140.846016
Rwneg12_96 in12 sn96 11140.846016
Rwneg12_97 in12 sn97 3183.098862
Rwneg12_98 in12 sn98 11140.846016
Rwneg12_99 in12 sn99 3183.098862
Rwneg12_100 in12 sn100 3183.098862
Rwneg13_1 in13 sn1 11140.846016
Rwneg13_2 in13 sn2 11140.846016
Rwneg13_3 in13 sn3 11140.846016
Rwneg13_4 in13 sn4 11140.846016
Rwneg13_5 in13 sn5 3183.098862
Rwneg13_6 in13 sn6 11140.846016
Rwneg13_7 in13 sn7 11140.846016
Rwneg13_8 in13 sn8 11140.846016
Rwneg13_9 in13 sn9 11140.846016
Rwneg13_10 in13 sn10 3183.098862
Rwneg13_11 in13 sn11 3183.098862
Rwneg13_12 in13 sn12 11140.846016
Rwneg13_13 in13 sn13 11140.846016
Rwneg13_14 in13 sn14 11140.846016
Rwneg13_15 in13 sn15 3183.098862
Rwneg13_16 in13 sn16 11140.846016
Rwneg13_17 in13 sn17 3183.098862
Rwneg13_18 in13 sn18 3183.098862
Rwneg13_19 in13 sn19 3183.098862
Rwneg13_20 in13 sn20 3183.098862
Rwneg13_21 in13 sn21 11140.846016
Rwneg13_22 in13 sn22 3183.098862
Rwneg13_23 in13 sn23 11140.846016
Rwneg13_24 in13 sn24 3183.098862
Rwneg13_25 in13 sn25 3183.098862
Rwneg13_26 in13 sn26 3183.098862
Rwneg13_27 in13 sn27 11140.846016
Rwneg13_28 in13 sn28 11140.846016
Rwneg13_29 in13 sn29 3183.098862
Rwneg13_30 in13 sn30 11140.846016
Rwneg13_31 in13 sn31 3183.098862
Rwneg13_32 in13 sn32 3183.098862
Rwneg13_33 in13 sn33 11140.846016
Rwneg13_34 in13 sn34 11140.846016
Rwneg13_35 in13 sn35 11140.846016
Rwneg13_36 in13 sn36 3183.098862
Rwneg13_37 in13 sn37 3183.098862
Rwneg13_38 in13 sn38 3183.098862
Rwneg13_39 in13 sn39 3183.098862
Rwneg13_40 in13 sn40 11140.846016
Rwneg13_41 in13 sn41 3183.098862
Rwneg13_42 in13 sn42 11140.846016
Rwneg13_43 in13 sn43 3183.098862
Rwneg13_44 in13 sn44 3183.098862
Rwneg13_45 in13 sn45 11140.846016
Rwneg13_46 in13 sn46 11140.846016
Rwneg13_47 in13 sn47 11140.846016
Rwneg13_48 in13 sn48 11140.846016
Rwneg13_49 in13 sn49 3183.098862
Rwneg13_50 in13 sn50 3183.098862
Rwneg13_51 in13 sn51 3183.098862
Rwneg13_52 in13 sn52 3183.098862
Rwneg13_53 in13 sn53 11140.846016
Rwneg13_54 in13 sn54 3183.098862
Rwneg13_55 in13 sn55 3183.098862
Rwneg13_56 in13 sn56 3183.098862
Rwneg13_57 in13 sn57 11140.846016
Rwneg13_58 in13 sn58 11140.846016
Rwneg13_59 in13 sn59 3183.098862
Rwneg13_60 in13 sn60 11140.846016
Rwneg13_61 in13 sn61 3183.098862
Rwneg13_62 in13 sn62 11140.846016
Rwneg13_63 in13 sn63 11140.846016
Rwneg13_64 in13 sn64 11140.846016
Rwneg13_65 in13 sn65 3183.098862
Rwneg13_66 in13 sn66 3183.098862
Rwneg13_67 in13 sn67 3183.098862
Rwneg13_68 in13 sn68 11140.846016
Rwneg13_69 in13 sn69 3183.098862
Rwneg13_70 in13 sn70 3183.098862
Rwneg13_71 in13 sn71 11140.846016
Rwneg13_72 in13 sn72 3183.098862
Rwneg13_73 in13 sn73 3183.098862
Rwneg13_74 in13 sn74 11140.846016
Rwneg13_75 in13 sn75 11140.846016
Rwneg13_76 in13 sn76 3183.098862
Rwneg13_77 in13 sn77 3183.098862
Rwneg13_78 in13 sn78 11140.846016
Rwneg13_79 in13 sn79 3183.098862
Rwneg13_80 in13 sn80 3183.098862
Rwneg13_81 in13 sn81 11140.846016
Rwneg13_82 in13 sn82 11140.846016
Rwneg13_83 in13 sn83 3183.098862
Rwneg13_84 in13 sn84 3183.098862
Rwneg13_85 in13 sn85 3183.098862
Rwneg13_86 in13 sn86 3183.098862
Rwneg13_87 in13 sn87 3183.098862
Rwneg13_88 in13 sn88 11140.846016
Rwneg13_89 in13 sn89 11140.846016
Rwneg13_90 in13 sn90 11140.846016
Rwneg13_91 in13 sn91 3183.098862
Rwneg13_92 in13 sn92 3183.098862
Rwneg13_93 in13 sn93 11140.846016
Rwneg13_94 in13 sn94 11140.846016
Rwneg13_95 in13 sn95 3183.098862
Rwneg13_96 in13 sn96 11140.846016
Rwneg13_97 in13 sn97 11140.846016
Rwneg13_98 in13 sn98 11140.846016
Rwneg13_99 in13 sn99 3183.098862
Rwneg13_100 in13 sn100 11140.846016
Rwneg14_1 in14 sn1 3183.098862
Rwneg14_2 in14 sn2 3183.098862
Rwneg14_3 in14 sn3 3183.098862
Rwneg14_4 in14 sn4 11140.846016
Rwneg14_5 in14 sn5 3183.098862
Rwneg14_6 in14 sn6 3183.098862
Rwneg14_7 in14 sn7 11140.846016
Rwneg14_8 in14 sn8 11140.846016
Rwneg14_9 in14 sn9 3183.098862
Rwneg14_10 in14 sn10 11140.846016
Rwneg14_11 in14 sn11 11140.846016
Rwneg14_12 in14 sn12 11140.846016
Rwneg14_13 in14 sn13 11140.846016
Rwneg14_14 in14 sn14 11140.846016
Rwneg14_15 in14 sn15 3183.098862
Rwneg14_16 in14 sn16 3183.098862
Rwneg14_17 in14 sn17 11140.846016
Rwneg14_18 in14 sn18 11140.846016
Rwneg14_19 in14 sn19 11140.846016
Rwneg14_20 in14 sn20 3183.098862
Rwneg14_21 in14 sn21 11140.846016
Rwneg14_22 in14 sn22 11140.846016
Rwneg14_23 in14 sn23 11140.846016
Rwneg14_24 in14 sn24 11140.846016
Rwneg14_25 in14 sn25 11140.846016
Rwneg14_26 in14 sn26 11140.846016
Rwneg14_27 in14 sn27 3183.098862
Rwneg14_28 in14 sn28 3183.098862
Rwneg14_29 in14 sn29 3183.098862
Rwneg14_30 in14 sn30 11140.846016
Rwneg14_31 in14 sn31 11140.846016
Rwneg14_32 in14 sn32 11140.846016
Rwneg14_33 in14 sn33 11140.846016
Rwneg14_34 in14 sn34 3183.098862
Rwneg14_35 in14 sn35 3183.098862
Rwneg14_36 in14 sn36 3183.098862
Rwneg14_37 in14 sn37 3183.098862
Rwneg14_38 in14 sn38 11140.846016
Rwneg14_39 in14 sn39 3183.098862
Rwneg14_40 in14 sn40 11140.846016
Rwneg14_41 in14 sn41 11140.846016
Rwneg14_42 in14 sn42 3183.098862
Rwneg14_43 in14 sn43 3183.098862
Rwneg14_44 in14 sn44 11140.846016
Rwneg14_45 in14 sn45 3183.098862
Rwneg14_46 in14 sn46 3183.098862
Rwneg14_47 in14 sn47 3183.098862
Rwneg14_48 in14 sn48 11140.846016
Rwneg14_49 in14 sn49 3183.098862
Rwneg14_50 in14 sn50 11140.846016
Rwneg14_51 in14 sn51 3183.098862
Rwneg14_52 in14 sn52 11140.846016
Rwneg14_53 in14 sn53 11140.846016
Rwneg14_54 in14 sn54 3183.098862
Rwneg14_55 in14 sn55 3183.098862
Rwneg14_56 in14 sn56 3183.098862
Rwneg14_57 in14 sn57 3183.098862
Rwneg14_58 in14 sn58 11140.846016
Rwneg14_59 in14 sn59 11140.846016
Rwneg14_60 in14 sn60 3183.098862
Rwneg14_61 in14 sn61 3183.098862
Rwneg14_62 in14 sn62 11140.846016
Rwneg14_63 in14 sn63 11140.846016
Rwneg14_64 in14 sn64 11140.846016
Rwneg14_65 in14 sn65 11140.846016
Rwneg14_66 in14 sn66 11140.846016
Rwneg14_67 in14 sn67 3183.098862
Rwneg14_68 in14 sn68 3183.098862
Rwneg14_69 in14 sn69 11140.846016
Rwneg14_70 in14 sn70 3183.098862
Rwneg14_71 in14 sn71 3183.098862
Rwneg14_72 in14 sn72 11140.846016
Rwneg14_73 in14 sn73 11140.846016
Rwneg14_74 in14 sn74 11140.846016
Rwneg14_75 in14 sn75 11140.846016
Rwneg14_76 in14 sn76 3183.098862
Rwneg14_77 in14 sn77 11140.846016
Rwneg14_78 in14 sn78 3183.098862
Rwneg14_79 in14 sn79 11140.846016
Rwneg14_80 in14 sn80 3183.098862
Rwneg14_81 in14 sn81 3183.098862
Rwneg14_82 in14 sn82 3183.098862
Rwneg14_83 in14 sn83 3183.098862
Rwneg14_84 in14 sn84 11140.846016
Rwneg14_85 in14 sn85 11140.846016
Rwneg14_86 in14 sn86 3183.098862
Rwneg14_87 in14 sn87 3183.098862
Rwneg14_88 in14 sn88 3183.098862
Rwneg14_89 in14 sn89 3183.098862
Rwneg14_90 in14 sn90 11140.846016
Rwneg14_91 in14 sn91 11140.846016
Rwneg14_92 in14 sn92 3183.098862
Rwneg14_93 in14 sn93 3183.098862
Rwneg14_94 in14 sn94 11140.846016
Rwneg14_95 in14 sn95 11140.846016
Rwneg14_96 in14 sn96 11140.846016
Rwneg14_97 in14 sn97 3183.098862
Rwneg14_98 in14 sn98 3183.098862
Rwneg14_99 in14 sn99 3183.098862
Rwneg14_100 in14 sn100 3183.098862
Rwneg15_1 in15 sn1 3183.098862
Rwneg15_2 in15 sn2 3183.098862
Rwneg15_3 in15 sn3 11140.846016
Rwneg15_4 in15 sn4 11140.846016
Rwneg15_5 in15 sn5 11140.846016
Rwneg15_6 in15 sn6 3183.098862
Rwneg15_7 in15 sn7 3183.098862
Rwneg15_8 in15 sn8 3183.098862
Rwneg15_9 in15 sn9 3183.098862
Rwneg15_10 in15 sn10 11140.846016
Rwneg15_11 in15 sn11 3183.098862
Rwneg15_12 in15 sn12 3183.098862
Rwneg15_13 in15 sn13 3183.098862
Rwneg15_14 in15 sn14 11140.846016
Rwneg15_15 in15 sn15 11140.846016
Rwneg15_16 in15 sn16 3183.098862
Rwneg15_17 in15 sn17 3183.098862
Rwneg15_18 in15 sn18 3183.098862
Rwneg15_19 in15 sn19 3183.098862
Rwneg15_20 in15 sn20 3183.098862
Rwneg15_21 in15 sn21 11140.846016
Rwneg15_22 in15 sn22 11140.846016
Rwneg15_23 in15 sn23 3183.098862
Rwneg15_24 in15 sn24 11140.846016
Rwneg15_25 in15 sn25 3183.098862
Rwneg15_26 in15 sn26 3183.098862
Rwneg15_27 in15 sn27 3183.098862
Rwneg15_28 in15 sn28 11140.846016
Rwneg15_29 in15 sn29 3183.098862
Rwneg15_30 in15 sn30 11140.846016
Rwneg15_31 in15 sn31 11140.846016
Rwneg15_32 in15 sn32 11140.846016
Rwneg15_33 in15 sn33 11140.846016
Rwneg15_34 in15 sn34 11140.846016
Rwneg15_35 in15 sn35 11140.846016
Rwneg15_36 in15 sn36 3183.098862
Rwneg15_37 in15 sn37 11140.846016
Rwneg15_38 in15 sn38 11140.846016
Rwneg15_39 in15 sn39 11140.846016
Rwneg15_40 in15 sn40 3183.098862
Rwneg15_41 in15 sn41 3183.098862
Rwneg15_42 in15 sn42 11140.846016
Rwneg15_43 in15 sn43 3183.098862
Rwneg15_44 in15 sn44 3183.098862
Rwneg15_45 in15 sn45 3183.098862
Rwneg15_46 in15 sn46 3183.098862
Rwneg15_47 in15 sn47 3183.098862
Rwneg15_48 in15 sn48 3183.098862
Rwneg15_49 in15 sn49 11140.846016
Rwneg15_50 in15 sn50 3183.098862
Rwneg15_51 in15 sn51 11140.846016
Rwneg15_52 in15 sn52 11140.846016
Rwneg15_53 in15 sn53 3183.098862
Rwneg15_54 in15 sn54 3183.098862
Rwneg15_55 in15 sn55 3183.098862
Rwneg15_56 in15 sn56 11140.846016
Rwneg15_57 in15 sn57 11140.846016
Rwneg15_58 in15 sn58 11140.846016
Rwneg15_59 in15 sn59 11140.846016
Rwneg15_60 in15 sn60 3183.098862
Rwneg15_61 in15 sn61 11140.846016
Rwneg15_62 in15 sn62 3183.098862
Rwneg15_63 in15 sn63 11140.846016
Rwneg15_64 in15 sn64 11140.846016
Rwneg15_65 in15 sn65 11140.846016
Rwneg15_66 in15 sn66 3183.098862
Rwneg15_67 in15 sn67 3183.098862
Rwneg15_68 in15 sn68 11140.846016
Rwneg15_69 in15 sn69 11140.846016
Rwneg15_70 in15 sn70 11140.846016
Rwneg15_71 in15 sn71 11140.846016
Rwneg15_72 in15 sn72 3183.098862
Rwneg15_73 in15 sn73 11140.846016
Rwneg15_74 in15 sn74 3183.098862
Rwneg15_75 in15 sn75 11140.846016
Rwneg15_76 in15 sn76 3183.098862
Rwneg15_77 in15 sn77 3183.098862
Rwneg15_78 in15 sn78 3183.098862
Rwneg15_79 in15 sn79 11140.846016
Rwneg15_80 in15 sn80 11140.846016
Rwneg15_81 in15 sn81 11140.846016
Rwneg15_82 in15 sn82 11140.846016
Rwneg15_83 in15 sn83 11140.846016
Rwneg15_84 in15 sn84 3183.098862
Rwneg15_85 in15 sn85 3183.098862
Rwneg15_86 in15 sn86 3183.098862
Rwneg15_87 in15 sn87 3183.098862
Rwneg15_88 in15 sn88 3183.098862
Rwneg15_89 in15 sn89 11140.846016
Rwneg15_90 in15 sn90 3183.098862
Rwneg15_91 in15 sn91 11140.846016
Rwneg15_92 in15 sn92 11140.846016
Rwneg15_93 in15 sn93 3183.098862
Rwneg15_94 in15 sn94 11140.846016
Rwneg15_95 in15 sn95 11140.846016
Rwneg15_96 in15 sn96 11140.846016
Rwneg15_97 in15 sn97 3183.098862
Rwneg15_98 in15 sn98 11140.846016
Rwneg15_99 in15 sn99 3183.098862
Rwneg15_100 in15 sn100 11140.846016
Rwneg16_1 in16 sn1 11140.846016
Rwneg16_2 in16 sn2 11140.846016
Rwneg16_3 in16 sn3 3183.098862
Rwneg16_4 in16 sn4 3183.098862
Rwneg16_5 in16 sn5 11140.846016
Rwneg16_6 in16 sn6 11140.846016
Rwneg16_7 in16 sn7 3183.098862
Rwneg16_8 in16 sn8 3183.098862
Rwneg16_9 in16 sn9 11140.846016
Rwneg16_10 in16 sn10 3183.098862
Rwneg16_11 in16 sn11 3183.098862
Rwneg16_12 in16 sn12 11140.846016
Rwneg16_13 in16 sn13 11140.846016
Rwneg16_14 in16 sn14 11140.846016
Rwneg16_15 in16 sn15 3183.098862
Rwneg16_16 in16 sn16 11140.846016
Rwneg16_17 in16 sn17 11140.846016
Rwneg16_18 in16 sn18 11140.846016
Rwneg16_19 in16 sn19 3183.098862
Rwneg16_20 in16 sn20 11140.846016
Rwneg16_21 in16 sn21 3183.098862
Rwneg16_22 in16 sn22 11140.846016
Rwneg16_23 in16 sn23 11140.846016
Rwneg16_24 in16 sn24 3183.098862
Rwneg16_25 in16 sn25 3183.098862
Rwneg16_26 in16 sn26 3183.098862
Rwneg16_27 in16 sn27 3183.098862
Rwneg16_28 in16 sn28 3183.098862
Rwneg16_29 in16 sn29 3183.098862
Rwneg16_30 in16 sn30 3183.098862
Rwneg16_31 in16 sn31 3183.098862
Rwneg16_32 in16 sn32 3183.098862
Rwneg16_33 in16 sn33 3183.098862
Rwneg16_34 in16 sn34 3183.098862
Rwneg16_35 in16 sn35 11140.846016
Rwneg16_36 in16 sn36 3183.098862
Rwneg16_37 in16 sn37 3183.098862
Rwneg16_38 in16 sn38 11140.846016
Rwneg16_39 in16 sn39 3183.098862
Rwneg16_40 in16 sn40 11140.846016
Rwneg16_41 in16 sn41 3183.098862
Rwneg16_42 in16 sn42 11140.846016
Rwneg16_43 in16 sn43 3183.098862
Rwneg16_44 in16 sn44 11140.846016
Rwneg16_45 in16 sn45 11140.846016
Rwneg16_46 in16 sn46 3183.098862
Rwneg16_47 in16 sn47 3183.098862
Rwneg16_48 in16 sn48 11140.846016
Rwneg16_49 in16 sn49 11140.846016
Rwneg16_50 in16 sn50 11140.846016
Rwneg16_51 in16 sn51 11140.846016
Rwneg16_52 in16 sn52 3183.098862
Rwneg16_53 in16 sn53 3183.098862
Rwneg16_54 in16 sn54 11140.846016
Rwneg16_55 in16 sn55 3183.098862
Rwneg16_56 in16 sn56 11140.846016
Rwneg16_57 in16 sn57 11140.846016
Rwneg16_58 in16 sn58 3183.098862
Rwneg16_59 in16 sn59 11140.846016
Rwneg16_60 in16 sn60 11140.846016
Rwneg16_61 in16 sn61 11140.846016
Rwneg16_62 in16 sn62 11140.846016
Rwneg16_63 in16 sn63 3183.098862
Rwneg16_64 in16 sn64 3183.098862
Rwneg16_65 in16 sn65 11140.846016
Rwneg16_66 in16 sn66 11140.846016
Rwneg16_67 in16 sn67 11140.846016
Rwneg16_68 in16 sn68 11140.846016
Rwneg16_69 in16 sn69 3183.098862
Rwneg16_70 in16 sn70 11140.846016
Rwneg16_71 in16 sn71 11140.846016
Rwneg16_72 in16 sn72 11140.846016
Rwneg16_73 in16 sn73 11140.846016
Rwneg16_74 in16 sn74 3183.098862
Rwneg16_75 in16 sn75 3183.098862
Rwneg16_76 in16 sn76 11140.846016
Rwneg16_77 in16 sn77 11140.846016
Rwneg16_78 in16 sn78 11140.846016
Rwneg16_79 in16 sn79 3183.098862
Rwneg16_80 in16 sn80 3183.098862
Rwneg16_81 in16 sn81 11140.846016
Rwneg16_82 in16 sn82 11140.846016
Rwneg16_83 in16 sn83 3183.098862
Rwneg16_84 in16 sn84 3183.098862
Rwneg16_85 in16 sn85 3183.098862
Rwneg16_86 in16 sn86 11140.846016
Rwneg16_87 in16 sn87 11140.846016
Rwneg16_88 in16 sn88 11140.846016
Rwneg16_89 in16 sn89 3183.098862
Rwneg16_90 in16 sn90 3183.098862
Rwneg16_91 in16 sn91 3183.098862
Rwneg16_92 in16 sn92 11140.846016
Rwneg16_93 in16 sn93 11140.846016
Rwneg16_94 in16 sn94 3183.098862
Rwneg16_95 in16 sn95 3183.098862
Rwneg16_96 in16 sn96 11140.846016
Rwneg16_97 in16 sn97 11140.846016
Rwneg16_98 in16 sn98 11140.846016
Rwneg16_99 in16 sn99 11140.846016
Rwneg16_100 in16 sn100 3183.098862
Rwneg17_1 in17 sn1 3183.098862
Rwneg17_2 in17 sn2 11140.846016
Rwneg17_3 in17 sn3 3183.098862
Rwneg17_4 in17 sn4 3183.098862
Rwneg17_5 in17 sn5 3183.098862
Rwneg17_6 in17 sn6 3183.098862
Rwneg17_7 in17 sn7 11140.846016
Rwneg17_8 in17 sn8 11140.846016
Rwneg17_9 in17 sn9 11140.846016
Rwneg17_10 in17 sn10 3183.098862
Rwneg17_11 in17 sn11 11140.846016
Rwneg17_12 in17 sn12 11140.846016
Rwneg17_13 in17 sn13 11140.846016
Rwneg17_14 in17 sn14 11140.846016
Rwneg17_15 in17 sn15 11140.846016
Rwneg17_16 in17 sn16 3183.098862
Rwneg17_17 in17 sn17 11140.846016
Rwneg17_18 in17 sn18 11140.846016
Rwneg17_19 in17 sn19 3183.098862
Rwneg17_20 in17 sn20 3183.098862
Rwneg17_21 in17 sn21 3183.098862
Rwneg17_22 in17 sn22 3183.098862
Rwneg17_23 in17 sn23 11140.846016
Rwneg17_24 in17 sn24 11140.846016
Rwneg17_25 in17 sn25 11140.846016
Rwneg17_26 in17 sn26 11140.846016
Rwneg17_27 in17 sn27 3183.098862
Rwneg17_28 in17 sn28 11140.846016
Rwneg17_29 in17 sn29 11140.846016
Rwneg17_30 in17 sn30 11140.846016
Rwneg17_31 in17 sn31 3183.098862
Rwneg17_32 in17 sn32 3183.098862
Rwneg17_33 in17 sn33 11140.846016
Rwneg17_34 in17 sn34 11140.846016
Rwneg17_35 in17 sn35 3183.098862
Rwneg17_36 in17 sn36 11140.846016
Rwneg17_37 in17 sn37 3183.098862
Rwneg17_38 in17 sn38 3183.098862
Rwneg17_39 in17 sn39 11140.846016
Rwneg17_40 in17 sn40 3183.098862
Rwneg17_41 in17 sn41 11140.846016
Rwneg17_42 in17 sn42 3183.098862
Rwneg17_43 in17 sn43 3183.098862
Rwneg17_44 in17 sn44 11140.846016
Rwneg17_45 in17 sn45 11140.846016
Rwneg17_46 in17 sn46 11140.846016
Rwneg17_47 in17 sn47 11140.846016
Rwneg17_48 in17 sn48 3183.098862
Rwneg17_49 in17 sn49 11140.846016
Rwneg17_50 in17 sn50 11140.846016
Rwneg17_51 in17 sn51 3183.098862
Rwneg17_52 in17 sn52 11140.846016
Rwneg17_53 in17 sn53 3183.098862
Rwneg17_54 in17 sn54 3183.098862
Rwneg17_55 in17 sn55 3183.098862
Rwneg17_56 in17 sn56 11140.846016
Rwneg17_57 in17 sn57 11140.846016
Rwneg17_58 in17 sn58 3183.098862
Rwneg17_59 in17 sn59 11140.846016
Rwneg17_60 in17 sn60 11140.846016
Rwneg17_61 in17 sn61 11140.846016
Rwneg17_62 in17 sn62 11140.846016
Rwneg17_63 in17 sn63 11140.846016
Rwneg17_64 in17 sn64 3183.098862
Rwneg17_65 in17 sn65 11140.846016
Rwneg17_66 in17 sn66 3183.098862
Rwneg17_67 in17 sn67 11140.846016
Rwneg17_68 in17 sn68 11140.846016
Rwneg17_69 in17 sn69 3183.098862
Rwneg17_70 in17 sn70 3183.098862
Rwneg17_71 in17 sn71 11140.846016
Rwneg17_72 in17 sn72 11140.846016
Rwneg17_73 in17 sn73 11140.846016
Rwneg17_74 in17 sn74 3183.098862
Rwneg17_75 in17 sn75 11140.846016
Rwneg17_76 in17 sn76 11140.846016
Rwneg17_77 in17 sn77 3183.098862
Rwneg17_78 in17 sn78 11140.846016
Rwneg17_79 in17 sn79 11140.846016
Rwneg17_80 in17 sn80 3183.098862
Rwneg17_81 in17 sn81 3183.098862
Rwneg17_82 in17 sn82 11140.846016
Rwneg17_83 in17 sn83 3183.098862
Rwneg17_84 in17 sn84 11140.846016
Rwneg17_85 in17 sn85 3183.098862
Rwneg17_86 in17 sn86 3183.098862
Rwneg17_87 in17 sn87 11140.846016
Rwneg17_88 in17 sn88 3183.098862
Rwneg17_89 in17 sn89 3183.098862
Rwneg17_90 in17 sn90 3183.098862
Rwneg17_91 in17 sn91 11140.846016
Rwneg17_92 in17 sn92 3183.098862
Rwneg17_93 in17 sn93 11140.846016
Rwneg17_94 in17 sn94 3183.098862
Rwneg17_95 in17 sn95 11140.846016
Rwneg17_96 in17 sn96 3183.098862
Rwneg17_97 in17 sn97 11140.846016
Rwneg17_98 in17 sn98 3183.098862
Rwneg17_99 in17 sn99 3183.098862
Rwneg17_100 in17 sn100 3183.098862
Rwneg18_1 in18 sn1 3183.098862
Rwneg18_2 in18 sn2 3183.098862
Rwneg18_3 in18 sn3 3183.098862
Rwneg18_4 in18 sn4 3183.098862
Rwneg18_5 in18 sn5 3183.098862
Rwneg18_6 in18 sn6 3183.098862
Rwneg18_7 in18 sn7 3183.098862
Rwneg18_8 in18 sn8 11140.846016
Rwneg18_9 in18 sn9 11140.846016
Rwneg18_10 in18 sn10 3183.098862
Rwneg18_11 in18 sn11 3183.098862
Rwneg18_12 in18 sn12 3183.098862
Rwneg18_13 in18 sn13 3183.098862
Rwneg18_14 in18 sn14 3183.098862
Rwneg18_15 in18 sn15 3183.098862
Rwneg18_16 in18 sn16 11140.846016
Rwneg18_17 in18 sn17 11140.846016
Rwneg18_18 in18 sn18 3183.098862
Rwneg18_19 in18 sn19 11140.846016
Rwneg18_20 in18 sn20 3183.098862
Rwneg18_21 in18 sn21 3183.098862
Rwneg18_22 in18 sn22 11140.846016
Rwneg18_23 in18 sn23 11140.846016
Rwneg18_24 in18 sn24 3183.098862
Rwneg18_25 in18 sn25 3183.098862
Rwneg18_26 in18 sn26 11140.846016
Rwneg18_27 in18 sn27 11140.846016
Rwneg18_28 in18 sn28 3183.098862
Rwneg18_29 in18 sn29 11140.846016
Rwneg18_30 in18 sn30 3183.098862
Rwneg18_31 in18 sn31 3183.098862
Rwneg18_32 in18 sn32 3183.098862
Rwneg18_33 in18 sn33 3183.098862
Rwneg18_34 in18 sn34 11140.846016
Rwneg18_35 in18 sn35 11140.846016
Rwneg18_36 in18 sn36 11140.846016
Rwneg18_37 in18 sn37 3183.098862
Rwneg18_38 in18 sn38 11140.846016
Rwneg18_39 in18 sn39 11140.846016
Rwneg18_40 in18 sn40 3183.098862
Rwneg18_41 in18 sn41 3183.098862
Rwneg18_42 in18 sn42 3183.098862
Rwneg18_43 in18 sn43 11140.846016
Rwneg18_44 in18 sn44 3183.098862
Rwneg18_45 in18 sn45 3183.098862
Rwneg18_46 in18 sn46 3183.098862
Rwneg18_47 in18 sn47 11140.846016
Rwneg18_48 in18 sn48 3183.098862
Rwneg18_49 in18 sn49 3183.098862
Rwneg18_50 in18 sn50 3183.098862
Rwneg18_51 in18 sn51 11140.846016
Rwneg18_52 in18 sn52 3183.098862
Rwneg18_53 in18 sn53 11140.846016
Rwneg18_54 in18 sn54 11140.846016
Rwneg18_55 in18 sn55 3183.098862
Rwneg18_56 in18 sn56 11140.846016
Rwneg18_57 in18 sn57 3183.098862
Rwneg18_58 in18 sn58 3183.098862
Rwneg18_59 in18 sn59 3183.098862
Rwneg18_60 in18 sn60 3183.098862
Rwneg18_61 in18 sn61 11140.846016
Rwneg18_62 in18 sn62 11140.846016
Rwneg18_63 in18 sn63 11140.846016
Rwneg18_64 in18 sn64 3183.098862
Rwneg18_65 in18 sn65 11140.846016
Rwneg18_66 in18 sn66 3183.098862
Rwneg18_67 in18 sn67 11140.846016
Rwneg18_68 in18 sn68 3183.098862
Rwneg18_69 in18 sn69 11140.846016
Rwneg18_70 in18 sn70 3183.098862
Rwneg18_71 in18 sn71 3183.098862
Rwneg18_72 in18 sn72 11140.846016
Rwneg18_73 in18 sn73 11140.846016
Rwneg18_74 in18 sn74 3183.098862
Rwneg18_75 in18 sn75 11140.846016
Rwneg18_76 in18 sn76 11140.846016
Rwneg18_77 in18 sn77 11140.846016
Rwneg18_78 in18 sn78 11140.846016
Rwneg18_79 in18 sn79 3183.098862
Rwneg18_80 in18 sn80 11140.846016
Rwneg18_81 in18 sn81 11140.846016
Rwneg18_82 in18 sn82 3183.098862
Rwneg18_83 in18 sn83 3183.098862
Rwneg18_84 in18 sn84 11140.846016
Rwneg18_85 in18 sn85 3183.098862
Rwneg18_86 in18 sn86 3183.098862
Rwneg18_87 in18 sn87 3183.098862
Rwneg18_88 in18 sn88 11140.846016
Rwneg18_89 in18 sn89 3183.098862
Rwneg18_90 in18 sn90 11140.846016
Rwneg18_91 in18 sn91 3183.098862
Rwneg18_92 in18 sn92 3183.098862
Rwneg18_93 in18 sn93 11140.846016
Rwneg18_94 in18 sn94 3183.098862
Rwneg18_95 in18 sn95 3183.098862
Rwneg18_96 in18 sn96 3183.098862
Rwneg18_97 in18 sn97 11140.846016
Rwneg18_98 in18 sn98 11140.846016
Rwneg18_99 in18 sn99 3183.098862
Rwneg18_100 in18 sn100 3183.098862
Rwneg19_1 in19 sn1 11140.846016
Rwneg19_2 in19 sn2 3183.098862
Rwneg19_3 in19 sn3 3183.098862
Rwneg19_4 in19 sn4 3183.098862
Rwneg19_5 in19 sn5 11140.846016
Rwneg19_6 in19 sn6 11140.846016
Rwneg19_7 in19 sn7 3183.098862
Rwneg19_8 in19 sn8 3183.098862
Rwneg19_9 in19 sn9 3183.098862
Rwneg19_10 in19 sn10 11140.846016
Rwneg19_11 in19 sn11 3183.098862
Rwneg19_12 in19 sn12 3183.098862
Rwneg19_13 in19 sn13 11140.846016
Rwneg19_14 in19 sn14 3183.098862
Rwneg19_15 in19 sn15 11140.846016
Rwneg19_16 in19 sn16 11140.846016
Rwneg19_17 in19 sn17 3183.098862
Rwneg19_18 in19 sn18 11140.846016
Rwneg19_19 in19 sn19 3183.098862
Rwneg19_20 in19 sn20 3183.098862
Rwneg19_21 in19 sn21 3183.098862
Rwneg19_22 in19 sn22 3183.098862
Rwneg19_23 in19 sn23 3183.098862
Rwneg19_24 in19 sn24 3183.098862
Rwneg19_25 in19 sn25 11140.846016
Rwneg19_26 in19 sn26 3183.098862
Rwneg19_27 in19 sn27 3183.098862
Rwneg19_28 in19 sn28 3183.098862
Rwneg19_29 in19 sn29 3183.098862
Rwneg19_30 in19 sn30 11140.846016
Rwneg19_31 in19 sn31 3183.098862
Rwneg19_32 in19 sn32 11140.846016
Rwneg19_33 in19 sn33 11140.846016
Rwneg19_34 in19 sn34 11140.846016
Rwneg19_35 in19 sn35 11140.846016
Rwneg19_36 in19 sn36 3183.098862
Rwneg19_37 in19 sn37 3183.098862
Rwneg19_38 in19 sn38 3183.098862
Rwneg19_39 in19 sn39 11140.846016
Rwneg19_40 in19 sn40 3183.098862
Rwneg19_41 in19 sn41 3183.098862
Rwneg19_42 in19 sn42 3183.098862
Rwneg19_43 in19 sn43 3183.098862
Rwneg19_44 in19 sn44 11140.846016
Rwneg19_45 in19 sn45 11140.846016
Rwneg19_46 in19 sn46 11140.846016
Rwneg19_47 in19 sn47 11140.846016
Rwneg19_48 in19 sn48 11140.846016
Rwneg19_49 in19 sn49 11140.846016
Rwneg19_50 in19 sn50 3183.098862
Rwneg19_51 in19 sn51 3183.098862
Rwneg19_52 in19 sn52 11140.846016
Rwneg19_53 in19 sn53 11140.846016
Rwneg19_54 in19 sn54 11140.846016
Rwneg19_55 in19 sn55 11140.846016
Rwneg19_56 in19 sn56 3183.098862
Rwneg19_57 in19 sn57 11140.846016
Rwneg19_58 in19 sn58 3183.098862
Rwneg19_59 in19 sn59 3183.098862
Rwneg19_60 in19 sn60 3183.098862
Rwneg19_61 in19 sn61 11140.846016
Rwneg19_62 in19 sn62 3183.098862
Rwneg19_63 in19 sn63 11140.846016
Rwneg19_64 in19 sn64 11140.846016
Rwneg19_65 in19 sn65 11140.846016
Rwneg19_66 in19 sn66 3183.098862
Rwneg19_67 in19 sn67 3183.098862
Rwneg19_68 in19 sn68 11140.846016
Rwneg19_69 in19 sn69 11140.846016
Rwneg19_70 in19 sn70 3183.098862
Rwneg19_71 in19 sn71 11140.846016
Rwneg19_72 in19 sn72 3183.098862
Rwneg19_73 in19 sn73 3183.098862
Rwneg19_74 in19 sn74 11140.846016
Rwneg19_75 in19 sn75 11140.846016
Rwneg19_76 in19 sn76 11140.846016
Rwneg19_77 in19 sn77 3183.098862
Rwneg19_78 in19 sn78 11140.846016
Rwneg19_79 in19 sn79 11140.846016
Rwneg19_80 in19 sn80 11140.846016
Rwneg19_81 in19 sn81 3183.098862
Rwneg19_82 in19 sn82 11140.846016
Rwneg19_83 in19 sn83 3183.098862
Rwneg19_84 in19 sn84 11140.846016
Rwneg19_85 in19 sn85 11140.846016
Rwneg19_86 in19 sn86 11140.846016
Rwneg19_87 in19 sn87 3183.098862
Rwneg19_88 in19 sn88 3183.098862
Rwneg19_89 in19 sn89 3183.098862
Rwneg19_90 in19 sn90 11140.846016
Rwneg19_91 in19 sn91 3183.098862
Rwneg19_92 in19 sn92 11140.846016
Rwneg19_93 in19 sn93 3183.098862
Rwneg19_94 in19 sn94 11140.846016
Rwneg19_95 in19 sn95 11140.846016
Rwneg19_96 in19 sn96 3183.098862
Rwneg19_97 in19 sn97 3183.098862
Rwneg19_98 in19 sn98 11140.846016
Rwneg19_99 in19 sn99 3183.098862
Rwneg19_100 in19 sn100 3183.098862
Rwneg20_1 in20 sn1 11140.846016
Rwneg20_2 in20 sn2 11140.846016
Rwneg20_3 in20 sn3 3183.098862
Rwneg20_4 in20 sn4 3183.098862
Rwneg20_5 in20 sn5 3183.098862
Rwneg20_6 in20 sn6 3183.098862
Rwneg20_7 in20 sn7 11140.846016
Rwneg20_8 in20 sn8 3183.098862
Rwneg20_9 in20 sn9 3183.098862
Rwneg20_10 in20 sn10 3183.098862
Rwneg20_11 in20 sn11 11140.846016
Rwneg20_12 in20 sn12 3183.098862
Rwneg20_13 in20 sn13 11140.846016
Rwneg20_14 in20 sn14 11140.846016
Rwneg20_15 in20 sn15 3183.098862
Rwneg20_16 in20 sn16 3183.098862
Rwneg20_17 in20 sn17 3183.098862
Rwneg20_18 in20 sn18 11140.846016
Rwneg20_19 in20 sn19 3183.098862
Rwneg20_20 in20 sn20 11140.846016
Rwneg20_21 in20 sn21 3183.098862
Rwneg20_22 in20 sn22 11140.846016
Rwneg20_23 in20 sn23 3183.098862
Rwneg20_24 in20 sn24 11140.846016
Rwneg20_25 in20 sn25 11140.846016
Rwneg20_26 in20 sn26 11140.846016
Rwneg20_27 in20 sn27 11140.846016
Rwneg20_28 in20 sn28 3183.098862
Rwneg20_29 in20 sn29 3183.098862
Rwneg20_30 in20 sn30 3183.098862
Rwneg20_31 in20 sn31 3183.098862
Rwneg20_32 in20 sn32 11140.846016
Rwneg20_33 in20 sn33 11140.846016
Rwneg20_34 in20 sn34 11140.846016
Rwneg20_35 in20 sn35 11140.846016
Rwneg20_36 in20 sn36 3183.098862
Rwneg20_37 in20 sn37 11140.846016
Rwneg20_38 in20 sn38 11140.846016
Rwneg20_39 in20 sn39 3183.098862
Rwneg20_40 in20 sn40 11140.846016
Rwneg20_41 in20 sn41 3183.098862
Rwneg20_42 in20 sn42 3183.098862
Rwneg20_43 in20 sn43 11140.846016
Rwneg20_44 in20 sn44 11140.846016
Rwneg20_45 in20 sn45 11140.846016
Rwneg20_46 in20 sn46 11140.846016
Rwneg20_47 in20 sn47 3183.098862
Rwneg20_48 in20 sn48 11140.846016
Rwneg20_49 in20 sn49 11140.846016
Rwneg20_50 in20 sn50 11140.846016
Rwneg20_51 in20 sn51 11140.846016
Rwneg20_52 in20 sn52 3183.098862
Rwneg20_53 in20 sn53 3183.098862
Rwneg20_54 in20 sn54 11140.846016
Rwneg20_55 in20 sn55 11140.846016
Rwneg20_56 in20 sn56 11140.846016
Rwneg20_57 in20 sn57 3183.098862
Rwneg20_58 in20 sn58 11140.846016
Rwneg20_59 in20 sn59 11140.846016
Rwneg20_60 in20 sn60 3183.098862
Rwneg20_61 in20 sn61 11140.846016
Rwneg20_62 in20 sn62 11140.846016
Rwneg20_63 in20 sn63 3183.098862
Rwneg20_64 in20 sn64 3183.098862
Rwneg20_65 in20 sn65 3183.098862
Rwneg20_66 in20 sn66 11140.846016
Rwneg20_67 in20 sn67 3183.098862
Rwneg20_68 in20 sn68 3183.098862
Rwneg20_69 in20 sn69 3183.098862
Rwneg20_70 in20 sn70 11140.846016
Rwneg20_71 in20 sn71 11140.846016
Rwneg20_72 in20 sn72 11140.846016
Rwneg20_73 in20 sn73 11140.846016
Rwneg20_74 in20 sn74 11140.846016
Rwneg20_75 in20 sn75 11140.846016
Rwneg20_76 in20 sn76 11140.846016
Rwneg20_77 in20 sn77 11140.846016
Rwneg20_78 in20 sn78 11140.846016
Rwneg20_79 in20 sn79 3183.098862
Rwneg20_80 in20 sn80 11140.846016
Rwneg20_81 in20 sn81 11140.846016
Rwneg20_82 in20 sn82 3183.098862
Rwneg20_83 in20 sn83 11140.846016
Rwneg20_84 in20 sn84 11140.846016
Rwneg20_85 in20 sn85 3183.098862
Rwneg20_86 in20 sn86 11140.846016
Rwneg20_87 in20 sn87 11140.846016
Rwneg20_88 in20 sn88 3183.098862
Rwneg20_89 in20 sn89 3183.098862
Rwneg20_90 in20 sn90 11140.846016
Rwneg20_91 in20 sn91 11140.846016
Rwneg20_92 in20 sn92 11140.846016
Rwneg20_93 in20 sn93 11140.846016
Rwneg20_94 in20 sn94 11140.846016
Rwneg20_95 in20 sn95 3183.098862
Rwneg20_96 in20 sn96 3183.098862
Rwneg20_97 in20 sn97 11140.846016
Rwneg20_98 in20 sn98 11140.846016
Rwneg20_99 in20 sn99 11140.846016
Rwneg20_100 in20 sn100 3183.098862
Rwneg21_1 in21 sn1 3183.098862
Rwneg21_2 in21 sn2 11140.846016
Rwneg21_3 in21 sn3 11140.846016
Rwneg21_4 in21 sn4 3183.098862
Rwneg21_5 in21 sn5 11140.846016
Rwneg21_6 in21 sn6 11140.846016
Rwneg21_7 in21 sn7 11140.846016
Rwneg21_8 in21 sn8 11140.846016
Rwneg21_9 in21 sn9 11140.846016
Rwneg21_10 in21 sn10 11140.846016
Rwneg21_11 in21 sn11 3183.098862
Rwneg21_12 in21 sn12 3183.098862
Rwneg21_13 in21 sn13 11140.846016
Rwneg21_14 in21 sn14 3183.098862
Rwneg21_15 in21 sn15 3183.098862
Rwneg21_16 in21 sn16 3183.098862
Rwneg21_17 in21 sn17 11140.846016
Rwneg21_18 in21 sn18 11140.846016
Rwneg21_19 in21 sn19 11140.846016
Rwneg21_20 in21 sn20 3183.098862
Rwneg21_21 in21 sn21 3183.098862
Rwneg21_22 in21 sn22 11140.846016
Rwneg21_23 in21 sn23 11140.846016
Rwneg21_24 in21 sn24 11140.846016
Rwneg21_25 in21 sn25 11140.846016
Rwneg21_26 in21 sn26 11140.846016
Rwneg21_27 in21 sn27 3183.098862
Rwneg21_28 in21 sn28 11140.846016
Rwneg21_29 in21 sn29 11140.846016
Rwneg21_30 in21 sn30 11140.846016
Rwneg21_31 in21 sn31 3183.098862
Rwneg21_32 in21 sn32 3183.098862
Rwneg21_33 in21 sn33 3183.098862
Rwneg21_34 in21 sn34 11140.846016
Rwneg21_35 in21 sn35 11140.846016
Rwneg21_36 in21 sn36 11140.846016
Rwneg21_37 in21 sn37 11140.846016
Rwneg21_38 in21 sn38 11140.846016
Rwneg21_39 in21 sn39 11140.846016
Rwneg21_40 in21 sn40 11140.846016
Rwneg21_41 in21 sn41 3183.098862
Rwneg21_42 in21 sn42 11140.846016
Rwneg21_43 in21 sn43 3183.098862
Rwneg21_44 in21 sn44 11140.846016
Rwneg21_45 in21 sn45 3183.098862
Rwneg21_46 in21 sn46 3183.098862
Rwneg21_47 in21 sn47 3183.098862
Rwneg21_48 in21 sn48 11140.846016
Rwneg21_49 in21 sn49 3183.098862
Rwneg21_50 in21 sn50 11140.846016
Rwneg21_51 in21 sn51 11140.846016
Rwneg21_52 in21 sn52 3183.098862
Rwneg21_53 in21 sn53 3183.098862
Rwneg21_54 in21 sn54 3183.098862
Rwneg21_55 in21 sn55 11140.846016
Rwneg21_56 in21 sn56 11140.846016
Rwneg21_57 in21 sn57 3183.098862
Rwneg21_58 in21 sn58 3183.098862
Rwneg21_59 in21 sn59 3183.098862
Rwneg21_60 in21 sn60 3183.098862
Rwneg21_61 in21 sn61 11140.846016
Rwneg21_62 in21 sn62 11140.846016
Rwneg21_63 in21 sn63 11140.846016
Rwneg21_64 in21 sn64 11140.846016
Rwneg21_65 in21 sn65 3183.098862
Rwneg21_66 in21 sn66 11140.846016
Rwneg21_67 in21 sn67 11140.846016
Rwneg21_68 in21 sn68 11140.846016
Rwneg21_69 in21 sn69 11140.846016
Rwneg21_70 in21 sn70 11140.846016
Rwneg21_71 in21 sn71 3183.098862
Rwneg21_72 in21 sn72 11140.846016
Rwneg21_73 in21 sn73 11140.846016
Rwneg21_74 in21 sn74 11140.846016
Rwneg21_75 in21 sn75 11140.846016
Rwneg21_76 in21 sn76 3183.098862
Rwneg21_77 in21 sn77 11140.846016
Rwneg21_78 in21 sn78 11140.846016
Rwneg21_79 in21 sn79 3183.098862
Rwneg21_80 in21 sn80 3183.098862
Rwneg21_81 in21 sn81 11140.846016
Rwneg21_82 in21 sn82 11140.846016
Rwneg21_83 in21 sn83 11140.846016
Rwneg21_84 in21 sn84 3183.098862
Rwneg21_85 in21 sn85 11140.846016
Rwneg21_86 in21 sn86 3183.098862
Rwneg21_87 in21 sn87 11140.846016
Rwneg21_88 in21 sn88 11140.846016
Rwneg21_89 in21 sn89 11140.846016
Rwneg21_90 in21 sn90 3183.098862
Rwneg21_91 in21 sn91 3183.098862
Rwneg21_92 in21 sn92 11140.846016
Rwneg21_93 in21 sn93 11140.846016
Rwneg21_94 in21 sn94 11140.846016
Rwneg21_95 in21 sn95 11140.846016
Rwneg21_96 in21 sn96 3183.098862
Rwneg21_97 in21 sn97 3183.098862
Rwneg21_98 in21 sn98 11140.846016
Rwneg21_99 in21 sn99 11140.846016
Rwneg21_100 in21 sn100 3183.098862
Rwneg22_1 in22 sn1 11140.846016
Rwneg22_2 in22 sn2 3183.098862
Rwneg22_3 in22 sn3 11140.846016
Rwneg22_4 in22 sn4 11140.846016
Rwneg22_5 in22 sn5 11140.846016
Rwneg22_6 in22 sn6 3183.098862
Rwneg22_7 in22 sn7 3183.098862
Rwneg22_8 in22 sn8 11140.846016
Rwneg22_9 in22 sn9 11140.846016
Rwneg22_10 in22 sn10 11140.846016
Rwneg22_11 in22 sn11 3183.098862
Rwneg22_12 in22 sn12 3183.098862
Rwneg22_13 in22 sn13 3183.098862
Rwneg22_14 in22 sn14 11140.846016
Rwneg22_15 in22 sn15 11140.846016
Rwneg22_16 in22 sn16 3183.098862
Rwneg22_17 in22 sn17 11140.846016
Rwneg22_18 in22 sn18 3183.098862
Rwneg22_19 in22 sn19 11140.846016
Rwneg22_20 in22 sn20 3183.098862
Rwneg22_21 in22 sn21 3183.098862
Rwneg22_22 in22 sn22 3183.098862
Rwneg22_23 in22 sn23 11140.846016
Rwneg22_24 in22 sn24 11140.846016
Rwneg22_25 in22 sn25 11140.846016
Rwneg22_26 in22 sn26 11140.846016
Rwneg22_27 in22 sn27 11140.846016
Rwneg22_28 in22 sn28 3183.098862
Rwneg22_29 in22 sn29 11140.846016
Rwneg22_30 in22 sn30 11140.846016
Rwneg22_31 in22 sn31 3183.098862
Rwneg22_32 in22 sn32 3183.098862
Rwneg22_33 in22 sn33 11140.846016
Rwneg22_34 in22 sn34 3183.098862
Rwneg22_35 in22 sn35 3183.098862
Rwneg22_36 in22 sn36 11140.846016
Rwneg22_37 in22 sn37 11140.846016
Rwneg22_38 in22 sn38 3183.098862
Rwneg22_39 in22 sn39 11140.846016
Rwneg22_40 in22 sn40 11140.846016
Rwneg22_41 in22 sn41 11140.846016
Rwneg22_42 in22 sn42 11140.846016
Rwneg22_43 in22 sn43 3183.098862
Rwneg22_44 in22 sn44 11140.846016
Rwneg22_45 in22 sn45 11140.846016
Rwneg22_46 in22 sn46 3183.098862
Rwneg22_47 in22 sn47 3183.098862
Rwneg22_48 in22 sn48 3183.098862
Rwneg22_49 in22 sn49 3183.098862
Rwneg22_50 in22 sn50 11140.846016
Rwneg22_51 in22 sn51 3183.098862
Rwneg22_52 in22 sn52 3183.098862
Rwneg22_53 in22 sn53 3183.098862
Rwneg22_54 in22 sn54 11140.846016
Rwneg22_55 in22 sn55 3183.098862
Rwneg22_56 in22 sn56 11140.846016
Rwneg22_57 in22 sn57 3183.098862
Rwneg22_58 in22 sn58 11140.846016
Rwneg22_59 in22 sn59 3183.098862
Rwneg22_60 in22 sn60 3183.098862
Rwneg22_61 in22 sn61 3183.098862
Rwneg22_62 in22 sn62 11140.846016
Rwneg22_63 in22 sn63 11140.846016
Rwneg22_64 in22 sn64 3183.098862
Rwneg22_65 in22 sn65 11140.846016
Rwneg22_66 in22 sn66 3183.098862
Rwneg22_67 in22 sn67 3183.098862
Rwneg22_68 in22 sn68 11140.846016
Rwneg22_69 in22 sn69 3183.098862
Rwneg22_70 in22 sn70 3183.098862
Rwneg22_71 in22 sn71 11140.846016
Rwneg22_72 in22 sn72 3183.098862
Rwneg22_73 in22 sn73 3183.098862
Rwneg22_74 in22 sn74 11140.846016
Rwneg22_75 in22 sn75 3183.098862
Rwneg22_76 in22 sn76 3183.098862
Rwneg22_77 in22 sn77 11140.846016
Rwneg22_78 in22 sn78 3183.098862
Rwneg22_79 in22 sn79 3183.098862
Rwneg22_80 in22 sn80 11140.846016
Rwneg22_81 in22 sn81 11140.846016
Rwneg22_82 in22 sn82 11140.846016
Rwneg22_83 in22 sn83 3183.098862
Rwneg22_84 in22 sn84 3183.098862
Rwneg22_85 in22 sn85 3183.098862
Rwneg22_86 in22 sn86 11140.846016
Rwneg22_87 in22 sn87 11140.846016
Rwneg22_88 in22 sn88 11140.846016
Rwneg22_89 in22 sn89 3183.098862
Rwneg22_90 in22 sn90 3183.098862
Rwneg22_91 in22 sn91 11140.846016
Rwneg22_92 in22 sn92 11140.846016
Rwneg22_93 in22 sn93 11140.846016
Rwneg22_94 in22 sn94 3183.098862
Rwneg22_95 in22 sn95 11140.846016
Rwneg22_96 in22 sn96 11140.846016
Rwneg22_97 in22 sn97 11140.846016
Rwneg22_98 in22 sn98 11140.846016
Rwneg22_99 in22 sn99 11140.846016
Rwneg22_100 in22 sn100 11140.846016
Rwneg23_1 in23 sn1 3183.098862
Rwneg23_2 in23 sn2 3183.098862
Rwneg23_3 in23 sn3 3183.098862
Rwneg23_4 in23 sn4 3183.098862
Rwneg23_5 in23 sn5 3183.098862
Rwneg23_6 in23 sn6 11140.846016
Rwneg23_7 in23 sn7 11140.846016
Rwneg23_8 in23 sn8 3183.098862
Rwneg23_9 in23 sn9 3183.098862
Rwneg23_10 in23 sn10 3183.098862
Rwneg23_11 in23 sn11 11140.846016
Rwneg23_12 in23 sn12 11140.846016
Rwneg23_13 in23 sn13 3183.098862
Rwneg23_14 in23 sn14 3183.098862
Rwneg23_15 in23 sn15 11140.846016
Rwneg23_16 in23 sn16 11140.846016
Rwneg23_17 in23 sn17 11140.846016
Rwneg23_18 in23 sn18 3183.098862
Rwneg23_19 in23 sn19 3183.098862
Rwneg23_20 in23 sn20 11140.846016
Rwneg23_21 in23 sn21 11140.846016
Rwneg23_22 in23 sn22 11140.846016
Rwneg23_23 in23 sn23 3183.098862
Rwneg23_24 in23 sn24 3183.098862
Rwneg23_25 in23 sn25 3183.098862
Rwneg23_26 in23 sn26 3183.098862
Rwneg23_27 in23 sn27 11140.846016
Rwneg23_28 in23 sn28 3183.098862
Rwneg23_29 in23 sn29 11140.846016
Rwneg23_30 in23 sn30 11140.846016
Rwneg23_31 in23 sn31 3183.098862
Rwneg23_32 in23 sn32 3183.098862
Rwneg23_33 in23 sn33 11140.846016
Rwneg23_34 in23 sn34 3183.098862
Rwneg23_35 in23 sn35 11140.846016
Rwneg23_36 in23 sn36 11140.846016
Rwneg23_37 in23 sn37 11140.846016
Rwneg23_38 in23 sn38 3183.098862
Rwneg23_39 in23 sn39 3183.098862
Rwneg23_40 in23 sn40 3183.098862
Rwneg23_41 in23 sn41 11140.846016
Rwneg23_42 in23 sn42 3183.098862
Rwneg23_43 in23 sn43 3183.098862
Rwneg23_44 in23 sn44 11140.846016
Rwneg23_45 in23 sn45 3183.098862
Rwneg23_46 in23 sn46 11140.846016
Rwneg23_47 in23 sn47 3183.098862
Rwneg23_48 in23 sn48 3183.098862
Rwneg23_49 in23 sn49 3183.098862
Rwneg23_50 in23 sn50 3183.098862
Rwneg23_51 in23 sn51 11140.846016
Rwneg23_52 in23 sn52 3183.098862
Rwneg23_53 in23 sn53 3183.098862
Rwneg23_54 in23 sn54 11140.846016
Rwneg23_55 in23 sn55 3183.098862
Rwneg23_56 in23 sn56 3183.098862
Rwneg23_57 in23 sn57 3183.098862
Rwneg23_58 in23 sn58 3183.098862
Rwneg23_59 in23 sn59 11140.846016
Rwneg23_60 in23 sn60 11140.846016
Rwneg23_61 in23 sn61 11140.846016
Rwneg23_62 in23 sn62 11140.846016
Rwneg23_63 in23 sn63 3183.098862
Rwneg23_64 in23 sn64 3183.098862
Rwneg23_65 in23 sn65 11140.846016
Rwneg23_66 in23 sn66 11140.846016
Rwneg23_67 in23 sn67 11140.846016
Rwneg23_68 in23 sn68 11140.846016
Rwneg23_69 in23 sn69 3183.098862
Rwneg23_70 in23 sn70 11140.846016
Rwneg23_71 in23 sn71 11140.846016
Rwneg23_72 in23 sn72 3183.098862
Rwneg23_73 in23 sn73 11140.846016
Rwneg23_74 in23 sn74 3183.098862
Rwneg23_75 in23 sn75 3183.098862
Rwneg23_76 in23 sn76 11140.846016
Rwneg23_77 in23 sn77 11140.846016
Rwneg23_78 in23 sn78 11140.846016
Rwneg23_79 in23 sn79 3183.098862
Rwneg23_80 in23 sn80 11140.846016
Rwneg23_81 in23 sn81 3183.098862
Rwneg23_82 in23 sn82 3183.098862
Rwneg23_83 in23 sn83 3183.098862
Rwneg23_84 in23 sn84 3183.098862
Rwneg23_85 in23 sn85 3183.098862
Rwneg23_86 in23 sn86 11140.846016
Rwneg23_87 in23 sn87 3183.098862
Rwneg23_88 in23 sn88 3183.098862
Rwneg23_89 in23 sn89 3183.098862
Rwneg23_90 in23 sn90 11140.846016
Rwneg23_91 in23 sn91 3183.098862
Rwneg23_92 in23 sn92 11140.846016
Rwneg23_93 in23 sn93 3183.098862
Rwneg23_94 in23 sn94 3183.098862
Rwneg23_95 in23 sn95 11140.846016
Rwneg23_96 in23 sn96 3183.098862
Rwneg23_97 in23 sn97 3183.098862
Rwneg23_98 in23 sn98 3183.098862
Rwneg23_99 in23 sn99 11140.846016
Rwneg23_100 in23 sn100 11140.846016
Rwneg24_1 in24 sn1 3183.098862
Rwneg24_2 in24 sn2 11140.846016
Rwneg24_3 in24 sn3 3183.098862
Rwneg24_4 in24 sn4 3183.098862
Rwneg24_5 in24 sn5 3183.098862
Rwneg24_6 in24 sn6 3183.098862
Rwneg24_7 in24 sn7 11140.846016
Rwneg24_8 in24 sn8 3183.098862
Rwneg24_9 in24 sn9 3183.098862
Rwneg24_10 in24 sn10 11140.846016
Rwneg24_11 in24 sn11 3183.098862
Rwneg24_12 in24 sn12 3183.098862
Rwneg24_13 in24 sn13 3183.098862
Rwneg24_14 in24 sn14 3183.098862
Rwneg24_15 in24 sn15 11140.846016
Rwneg24_16 in24 sn16 3183.098862
Rwneg24_17 in24 sn17 3183.098862
Rwneg24_18 in24 sn18 11140.846016
Rwneg24_19 in24 sn19 11140.846016
Rwneg24_20 in24 sn20 3183.098862
Rwneg24_21 in24 sn21 11140.846016
Rwneg24_22 in24 sn22 3183.098862
Rwneg24_23 in24 sn23 3183.098862
Rwneg24_24 in24 sn24 11140.846016
Rwneg24_25 in24 sn25 3183.098862
Rwneg24_26 in24 sn26 11140.846016
Rwneg24_27 in24 sn27 11140.846016
Rwneg24_28 in24 sn28 3183.098862
Rwneg24_29 in24 sn29 3183.098862
Rwneg24_30 in24 sn30 3183.098862
Rwneg24_31 in24 sn31 3183.098862
Rwneg24_32 in24 sn32 11140.846016
Rwneg24_33 in24 sn33 11140.846016
Rwneg24_34 in24 sn34 3183.098862
Rwneg24_35 in24 sn35 11140.846016
Rwneg24_36 in24 sn36 3183.098862
Rwneg24_37 in24 sn37 11140.846016
Rwneg24_38 in24 sn38 3183.098862
Rwneg24_39 in24 sn39 3183.098862
Rwneg24_40 in24 sn40 11140.846016
Rwneg24_41 in24 sn41 3183.098862
Rwneg24_42 in24 sn42 3183.098862
Rwneg24_43 in24 sn43 11140.846016
Rwneg24_44 in24 sn44 3183.098862
Rwneg24_45 in24 sn45 11140.846016
Rwneg24_46 in24 sn46 11140.846016
Rwneg24_47 in24 sn47 3183.098862
Rwneg24_48 in24 sn48 3183.098862
Rwneg24_49 in24 sn49 3183.098862
Rwneg24_50 in24 sn50 3183.098862
Rwneg24_51 in24 sn51 11140.846016
Rwneg24_52 in24 sn52 11140.846016
Rwneg24_53 in24 sn53 3183.098862
Rwneg24_54 in24 sn54 11140.846016
Rwneg24_55 in24 sn55 11140.846016
Rwneg24_56 in24 sn56 11140.846016
Rwneg24_57 in24 sn57 3183.098862
Rwneg24_58 in24 sn58 11140.846016
Rwneg24_59 in24 sn59 3183.098862
Rwneg24_60 in24 sn60 11140.846016
Rwneg24_61 in24 sn61 11140.846016
Rwneg24_62 in24 sn62 11140.846016
Rwneg24_63 in24 sn63 3183.098862
Rwneg24_64 in24 sn64 3183.098862
Rwneg24_65 in24 sn65 3183.098862
Rwneg24_66 in24 sn66 11140.846016
Rwneg24_67 in24 sn67 11140.846016
Rwneg24_68 in24 sn68 11140.846016
Rwneg24_69 in24 sn69 3183.098862
Rwneg24_70 in24 sn70 11140.846016
Rwneg24_71 in24 sn71 11140.846016
Rwneg24_72 in24 sn72 3183.098862
Rwneg24_73 in24 sn73 3183.098862
Rwneg24_74 in24 sn74 3183.098862
Rwneg24_75 in24 sn75 11140.846016
Rwneg24_76 in24 sn76 3183.098862
Rwneg24_77 in24 sn77 11140.846016
Rwneg24_78 in24 sn78 11140.846016
Rwneg24_79 in24 sn79 3183.098862
Rwneg24_80 in24 sn80 11140.846016
Rwneg24_81 in24 sn81 11140.846016
Rwneg24_82 in24 sn82 11140.846016
Rwneg24_83 in24 sn83 11140.846016
Rwneg24_84 in24 sn84 3183.098862
Rwneg24_85 in24 sn85 3183.098862
Rwneg24_86 in24 sn86 11140.846016
Rwneg24_87 in24 sn87 11140.846016
Rwneg24_88 in24 sn88 11140.846016
Rwneg24_89 in24 sn89 11140.846016
Rwneg24_90 in24 sn90 3183.098862
Rwneg24_91 in24 sn91 3183.098862
Rwneg24_92 in24 sn92 11140.846016
Rwneg24_93 in24 sn93 11140.846016
Rwneg24_94 in24 sn94 3183.098862
Rwneg24_95 in24 sn95 3183.098862
Rwneg24_96 in24 sn96 3183.098862
Rwneg24_97 in24 sn97 11140.846016
Rwneg24_98 in24 sn98 11140.846016
Rwneg24_99 in24 sn99 11140.846016
Rwneg24_100 in24 sn100 11140.846016
Rwneg25_1 in25 sn1 11140.846016
Rwneg25_2 in25 sn2 11140.846016
Rwneg25_3 in25 sn3 11140.846016
Rwneg25_4 in25 sn4 11140.846016
Rwneg25_5 in25 sn5 11140.846016
Rwneg25_6 in25 sn6 3183.098862
Rwneg25_7 in25 sn7 11140.846016
Rwneg25_8 in25 sn8 3183.098862
Rwneg25_9 in25 sn9 3183.098862
Rwneg25_10 in25 sn10 11140.846016
Rwneg25_11 in25 sn11 3183.098862
Rwneg25_12 in25 sn12 3183.098862
Rwneg25_13 in25 sn13 11140.846016
Rwneg25_14 in25 sn14 3183.098862
Rwneg25_15 in25 sn15 11140.846016
Rwneg25_16 in25 sn16 3183.098862
Rwneg25_17 in25 sn17 3183.098862
Rwneg25_18 in25 sn18 11140.846016
Rwneg25_19 in25 sn19 11140.846016
Rwneg25_20 in25 sn20 11140.846016
Rwneg25_21 in25 sn21 3183.098862
Rwneg25_22 in25 sn22 11140.846016
Rwneg25_23 in25 sn23 11140.846016
Rwneg25_24 in25 sn24 3183.098862
Rwneg25_25 in25 sn25 11140.846016
Rwneg25_26 in25 sn26 11140.846016
Rwneg25_27 in25 sn27 3183.098862
Rwneg25_28 in25 sn28 3183.098862
Rwneg25_29 in25 sn29 11140.846016
Rwneg25_30 in25 sn30 11140.846016
Rwneg25_31 in25 sn31 11140.846016
Rwneg25_32 in25 sn32 3183.098862
Rwneg25_33 in25 sn33 11140.846016
Rwneg25_34 in25 sn34 3183.098862
Rwneg25_35 in25 sn35 11140.846016
Rwneg25_36 in25 sn36 11140.846016
Rwneg25_37 in25 sn37 11140.846016
Rwneg25_38 in25 sn38 3183.098862
Rwneg25_39 in25 sn39 11140.846016
Rwneg25_40 in25 sn40 11140.846016
Rwneg25_41 in25 sn41 11140.846016
Rwneg25_42 in25 sn42 3183.098862
Rwneg25_43 in25 sn43 3183.098862
Rwneg25_44 in25 sn44 11140.846016
Rwneg25_45 in25 sn45 3183.098862
Rwneg25_46 in25 sn46 3183.098862
Rwneg25_47 in25 sn47 11140.846016
Rwneg25_48 in25 sn48 11140.846016
Rwneg25_49 in25 sn49 3183.098862
Rwneg25_50 in25 sn50 3183.098862
Rwneg25_51 in25 sn51 11140.846016
Rwneg25_52 in25 sn52 11140.846016
Rwneg25_53 in25 sn53 11140.846016
Rwneg25_54 in25 sn54 11140.846016
Rwneg25_55 in25 sn55 11140.846016
Rwneg25_56 in25 sn56 11140.846016
Rwneg25_57 in25 sn57 3183.098862
Rwneg25_58 in25 sn58 11140.846016
Rwneg25_59 in25 sn59 3183.098862
Rwneg25_60 in25 sn60 3183.098862
Rwneg25_61 in25 sn61 11140.846016
Rwneg25_62 in25 sn62 11140.846016
Rwneg25_63 in25 sn63 11140.846016
Rwneg25_64 in25 sn64 11140.846016
Rwneg25_65 in25 sn65 11140.846016
Rwneg25_66 in25 sn66 3183.098862
Rwneg25_67 in25 sn67 11140.846016
Rwneg25_68 in25 sn68 11140.846016
Rwneg25_69 in25 sn69 11140.846016
Rwneg25_70 in25 sn70 11140.846016
Rwneg25_71 in25 sn71 11140.846016
Rwneg25_72 in25 sn72 11140.846016
Rwneg25_73 in25 sn73 11140.846016
Rwneg25_74 in25 sn74 11140.846016
Rwneg25_75 in25 sn75 3183.098862
Rwneg25_76 in25 sn76 3183.098862
Rwneg25_77 in25 sn77 3183.098862
Rwneg25_78 in25 sn78 3183.098862
Rwneg25_79 in25 sn79 3183.098862
Rwneg25_80 in25 sn80 11140.846016
Rwneg25_81 in25 sn81 11140.846016
Rwneg25_82 in25 sn82 3183.098862
Rwneg25_83 in25 sn83 11140.846016
Rwneg25_84 in25 sn84 11140.846016
Rwneg25_85 in25 sn85 3183.098862
Rwneg25_86 in25 sn86 3183.098862
Rwneg25_87 in25 sn87 11140.846016
Rwneg25_88 in25 sn88 11140.846016
Rwneg25_89 in25 sn89 11140.846016
Rwneg25_90 in25 sn90 11140.846016
Rwneg25_91 in25 sn91 3183.098862
Rwneg25_92 in25 sn92 3183.098862
Rwneg25_93 in25 sn93 11140.846016
Rwneg25_94 in25 sn94 3183.098862
Rwneg25_95 in25 sn95 3183.098862
Rwneg25_96 in25 sn96 3183.098862
Rwneg25_97 in25 sn97 11140.846016
Rwneg25_98 in25 sn98 3183.098862
Rwneg25_99 in25 sn99 11140.846016
Rwneg25_100 in25 sn100 11140.846016
Rwneg26_1 in26 sn1 11140.846016
Rwneg26_2 in26 sn2 3183.098862
Rwneg26_3 in26 sn3 11140.846016
Rwneg26_4 in26 sn4 11140.846016
Rwneg26_5 in26 sn5 3183.098862
Rwneg26_6 in26 sn6 11140.846016
Rwneg26_7 in26 sn7 3183.098862
Rwneg26_8 in26 sn8 3183.098862
Rwneg26_9 in26 sn9 3183.098862
Rwneg26_10 in26 sn10 3183.098862
Rwneg26_11 in26 sn11 11140.846016
Rwneg26_12 in26 sn12 3183.098862
Rwneg26_13 in26 sn13 11140.846016
Rwneg26_14 in26 sn14 3183.098862
Rwneg26_15 in26 sn15 11140.846016
Rwneg26_16 in26 sn16 11140.846016
Rwneg26_17 in26 sn17 11140.846016
Rwneg26_18 in26 sn18 11140.846016
Rwneg26_19 in26 sn19 11140.846016
Rwneg26_20 in26 sn20 11140.846016
Rwneg26_21 in26 sn21 3183.098862
Rwneg26_22 in26 sn22 11140.846016
Rwneg26_23 in26 sn23 11140.846016
Rwneg26_24 in26 sn24 3183.098862
Rwneg26_25 in26 sn25 3183.098862
Rwneg26_26 in26 sn26 3183.098862
Rwneg26_27 in26 sn27 11140.846016
Rwneg26_28 in26 sn28 11140.846016
Rwneg26_29 in26 sn29 11140.846016
Rwneg26_30 in26 sn30 3183.098862
Rwneg26_31 in26 sn31 11140.846016
Rwneg26_32 in26 sn32 11140.846016
Rwneg26_33 in26 sn33 11140.846016
Rwneg26_34 in26 sn34 3183.098862
Rwneg26_35 in26 sn35 11140.846016
Rwneg26_36 in26 sn36 11140.846016
Rwneg26_37 in26 sn37 3183.098862
Rwneg26_38 in26 sn38 3183.098862
Rwneg26_39 in26 sn39 3183.098862
Rwneg26_40 in26 sn40 3183.098862
Rwneg26_41 in26 sn41 11140.846016
Rwneg26_42 in26 sn42 3183.098862
Rwneg26_43 in26 sn43 3183.098862
Rwneg26_44 in26 sn44 3183.098862
Rwneg26_45 in26 sn45 11140.846016
Rwneg26_46 in26 sn46 11140.846016
Rwneg26_47 in26 sn47 11140.846016
Rwneg26_48 in26 sn48 3183.098862
Rwneg26_49 in26 sn49 11140.846016
Rwneg26_50 in26 sn50 11140.846016
Rwneg26_51 in26 sn51 11140.846016
Rwneg26_52 in26 sn52 11140.846016
Rwneg26_53 in26 sn53 3183.098862
Rwneg26_54 in26 sn54 11140.846016
Rwneg26_55 in26 sn55 11140.846016
Rwneg26_56 in26 sn56 3183.098862
Rwneg26_57 in26 sn57 3183.098862
Rwneg26_58 in26 sn58 11140.846016
Rwneg26_59 in26 sn59 3183.098862
Rwneg26_60 in26 sn60 11140.846016
Rwneg26_61 in26 sn61 11140.846016
Rwneg26_62 in26 sn62 3183.098862
Rwneg26_63 in26 sn63 11140.846016
Rwneg26_64 in26 sn64 3183.098862
Rwneg26_65 in26 sn65 11140.846016
Rwneg26_66 in26 sn66 3183.098862
Rwneg26_67 in26 sn67 3183.098862
Rwneg26_68 in26 sn68 3183.098862
Rwneg26_69 in26 sn69 11140.846016
Rwneg26_70 in26 sn70 3183.098862
Rwneg26_71 in26 sn71 11140.846016
Rwneg26_72 in26 sn72 11140.846016
Rwneg26_73 in26 sn73 3183.098862
Rwneg26_74 in26 sn74 11140.846016
Rwneg26_75 in26 sn75 11140.846016
Rwneg26_76 in26 sn76 3183.098862
Rwneg26_77 in26 sn77 11140.846016
Rwneg26_78 in26 sn78 11140.846016
Rwneg26_79 in26 sn79 11140.846016
Rwneg26_80 in26 sn80 3183.098862
Rwneg26_81 in26 sn81 11140.846016
Rwneg26_82 in26 sn82 11140.846016
Rwneg26_83 in26 sn83 3183.098862
Rwneg26_84 in26 sn84 11140.846016
Rwneg26_85 in26 sn85 3183.098862
Rwneg26_86 in26 sn86 11140.846016
Rwneg26_87 in26 sn87 11140.846016
Rwneg26_88 in26 sn88 3183.098862
Rwneg26_89 in26 sn89 11140.846016
Rwneg26_90 in26 sn90 3183.098862
Rwneg26_91 in26 sn91 3183.098862
Rwneg26_92 in26 sn92 11140.846016
Rwneg26_93 in26 sn93 11140.846016
Rwneg26_94 in26 sn94 3183.098862
Rwneg26_95 in26 sn95 11140.846016
Rwneg26_96 in26 sn96 3183.098862
Rwneg26_97 in26 sn97 11140.846016
Rwneg26_98 in26 sn98 3183.098862
Rwneg26_99 in26 sn99 3183.098862
Rwneg26_100 in26 sn100 11140.846016
Rwneg27_1 in27 sn1 11140.846016
Rwneg27_2 in27 sn2 3183.098862
Rwneg27_3 in27 sn3 11140.846016
Rwneg27_4 in27 sn4 11140.846016
Rwneg27_5 in27 sn5 3183.098862
Rwneg27_6 in27 sn6 11140.846016
Rwneg27_7 in27 sn7 11140.846016
Rwneg27_8 in27 sn8 3183.098862
Rwneg27_9 in27 sn9 11140.846016
Rwneg27_10 in27 sn10 3183.098862
Rwneg27_11 in27 sn11 3183.098862
Rwneg27_12 in27 sn12 3183.098862
Rwneg27_13 in27 sn13 3183.098862
Rwneg27_14 in27 sn14 11140.846016
Rwneg27_15 in27 sn15 3183.098862
Rwneg27_16 in27 sn16 3183.098862
Rwneg27_17 in27 sn17 11140.846016
Rwneg27_18 in27 sn18 3183.098862
Rwneg27_19 in27 sn19 11140.846016
Rwneg27_20 in27 sn20 11140.846016
Rwneg27_21 in27 sn21 3183.098862
Rwneg27_22 in27 sn22 11140.846016
Rwneg27_23 in27 sn23 11140.846016
Rwneg27_24 in27 sn24 3183.098862
Rwneg27_25 in27 sn25 11140.846016
Rwneg27_26 in27 sn26 11140.846016
Rwneg27_27 in27 sn27 11140.846016
Rwneg27_28 in27 sn28 11140.846016
Rwneg27_29 in27 sn29 3183.098862
Rwneg27_30 in27 sn30 11140.846016
Rwneg27_31 in27 sn31 3183.098862
Rwneg27_32 in27 sn32 3183.098862
Rwneg27_33 in27 sn33 3183.098862
Rwneg27_34 in27 sn34 3183.098862
Rwneg27_35 in27 sn35 11140.846016
Rwneg27_36 in27 sn36 11140.846016
Rwneg27_37 in27 sn37 3183.098862
Rwneg27_38 in27 sn38 11140.846016
Rwneg27_39 in27 sn39 11140.846016
Rwneg27_40 in27 sn40 11140.846016
Rwneg27_41 in27 sn41 3183.098862
Rwneg27_42 in27 sn42 11140.846016
Rwneg27_43 in27 sn43 3183.098862
Rwneg27_44 in27 sn44 11140.846016
Rwneg27_45 in27 sn45 11140.846016
Rwneg27_46 in27 sn46 11140.846016
Rwneg27_47 in27 sn47 11140.846016
Rwneg27_48 in27 sn48 11140.846016
Rwneg27_49 in27 sn49 3183.098862
Rwneg27_50 in27 sn50 11140.846016
Rwneg27_51 in27 sn51 11140.846016
Rwneg27_52 in27 sn52 11140.846016
Rwneg27_53 in27 sn53 11140.846016
Rwneg27_54 in27 sn54 3183.098862
Rwneg27_55 in27 sn55 3183.098862
Rwneg27_56 in27 sn56 11140.846016
Rwneg27_57 in27 sn57 3183.098862
Rwneg27_58 in27 sn58 3183.098862
Rwneg27_59 in27 sn59 3183.098862
Rwneg27_60 in27 sn60 3183.098862
Rwneg27_61 in27 sn61 11140.846016
Rwneg27_62 in27 sn62 11140.846016
Rwneg27_63 in27 sn63 11140.846016
Rwneg27_64 in27 sn64 11140.846016
Rwneg27_65 in27 sn65 11140.846016
Rwneg27_66 in27 sn66 3183.098862
Rwneg27_67 in27 sn67 11140.846016
Rwneg27_68 in27 sn68 11140.846016
Rwneg27_69 in27 sn69 11140.846016
Rwneg27_70 in27 sn70 11140.846016
Rwneg27_71 in27 sn71 11140.846016
Rwneg27_72 in27 sn72 11140.846016
Rwneg27_73 in27 sn73 3183.098862
Rwneg27_74 in27 sn74 11140.846016
Rwneg27_75 in27 sn75 3183.098862
Rwneg27_76 in27 sn76 11140.846016
Rwneg27_77 in27 sn77 3183.098862
Rwneg27_78 in27 sn78 11140.846016
Rwneg27_79 in27 sn79 3183.098862
Rwneg27_80 in27 sn80 11140.846016
Rwneg27_81 in27 sn81 11140.846016
Rwneg27_82 in27 sn82 3183.098862
Rwneg27_83 in27 sn83 11140.846016
Rwneg27_84 in27 sn84 3183.098862
Rwneg27_85 in27 sn85 11140.846016
Rwneg27_86 in27 sn86 11140.846016
Rwneg27_87 in27 sn87 3183.098862
Rwneg27_88 in27 sn88 3183.098862
Rwneg27_89 in27 sn89 11140.846016
Rwneg27_90 in27 sn90 11140.846016
Rwneg27_91 in27 sn91 3183.098862
Rwneg27_92 in27 sn92 3183.098862
Rwneg27_93 in27 sn93 3183.098862
Rwneg27_94 in27 sn94 3183.098862
Rwneg27_95 in27 sn95 11140.846016
Rwneg27_96 in27 sn96 11140.846016
Rwneg27_97 in27 sn97 3183.098862
Rwneg27_98 in27 sn98 11140.846016
Rwneg27_99 in27 sn99 11140.846016
Rwneg27_100 in27 sn100 3183.098862
Rwneg28_1 in28 sn1 3183.098862
Rwneg28_2 in28 sn2 3183.098862
Rwneg28_3 in28 sn3 11140.846016
Rwneg28_4 in28 sn4 11140.846016
Rwneg28_5 in28 sn5 11140.846016
Rwneg28_6 in28 sn6 3183.098862
Rwneg28_7 in28 sn7 3183.098862
Rwneg28_8 in28 sn8 11140.846016
Rwneg28_9 in28 sn9 3183.098862
Rwneg28_10 in28 sn10 3183.098862
Rwneg28_11 in28 sn11 3183.098862
Rwneg28_12 in28 sn12 3183.098862
Rwneg28_13 in28 sn13 3183.098862
Rwneg28_14 in28 sn14 11140.846016
Rwneg28_15 in28 sn15 3183.098862
Rwneg28_16 in28 sn16 3183.098862
Rwneg28_17 in28 sn17 11140.846016
Rwneg28_18 in28 sn18 11140.846016
Rwneg28_19 in28 sn19 11140.846016
Rwneg28_20 in28 sn20 3183.098862
Rwneg28_21 in28 sn21 3183.098862
Rwneg28_22 in28 sn22 3183.098862
Rwneg28_23 in28 sn23 3183.098862
Rwneg28_24 in28 sn24 3183.098862
Rwneg28_25 in28 sn25 11140.846016
Rwneg28_26 in28 sn26 11140.846016
Rwneg28_27 in28 sn27 11140.846016
Rwneg28_28 in28 sn28 11140.846016
Rwneg28_29 in28 sn29 3183.098862
Rwneg28_30 in28 sn30 11140.846016
Rwneg28_31 in28 sn31 11140.846016
Rwneg28_32 in28 sn32 11140.846016
Rwneg28_33 in28 sn33 3183.098862
Rwneg28_34 in28 sn34 11140.846016
Rwneg28_35 in28 sn35 11140.846016
Rwneg28_36 in28 sn36 11140.846016
Rwneg28_37 in28 sn37 11140.846016
Rwneg28_38 in28 sn38 3183.098862
Rwneg28_39 in28 sn39 11140.846016
Rwneg28_40 in28 sn40 3183.098862
Rwneg28_41 in28 sn41 11140.846016
Rwneg28_42 in28 sn42 11140.846016
Rwneg28_43 in28 sn43 11140.846016
Rwneg28_44 in28 sn44 3183.098862
Rwneg28_45 in28 sn45 3183.098862
Rwneg28_46 in28 sn46 11140.846016
Rwneg28_47 in28 sn47 3183.098862
Rwneg28_48 in28 sn48 11140.846016
Rwneg28_49 in28 sn49 11140.846016
Rwneg28_50 in28 sn50 11140.846016
Rwneg28_51 in28 sn51 3183.098862
Rwneg28_52 in28 sn52 11140.846016
Rwneg28_53 in28 sn53 11140.846016
Rwneg28_54 in28 sn54 3183.098862
Rwneg28_55 in28 sn55 3183.098862
Rwneg28_56 in28 sn56 3183.098862
Rwneg28_57 in28 sn57 11140.846016
Rwneg28_58 in28 sn58 3183.098862
Rwneg28_59 in28 sn59 3183.098862
Rwneg28_60 in28 sn60 11140.846016
Rwneg28_61 in28 sn61 11140.846016
Rwneg28_62 in28 sn62 11140.846016
Rwneg28_63 in28 sn63 3183.098862
Rwneg28_64 in28 sn64 11140.846016
Rwneg28_65 in28 sn65 11140.846016
Rwneg28_66 in28 sn66 3183.098862
Rwneg28_67 in28 sn67 11140.846016
Rwneg28_68 in28 sn68 11140.846016
Rwneg28_69 in28 sn69 3183.098862
Rwneg28_70 in28 sn70 11140.846016
Rwneg28_71 in28 sn71 3183.098862
Rwneg28_72 in28 sn72 11140.846016
Rwneg28_73 in28 sn73 3183.098862
Rwneg28_74 in28 sn74 3183.098862
Rwneg28_75 in28 sn75 3183.098862
Rwneg28_76 in28 sn76 11140.846016
Rwneg28_77 in28 sn77 11140.846016
Rwneg28_78 in28 sn78 11140.846016
Rwneg28_79 in28 sn79 3183.098862
Rwneg28_80 in28 sn80 11140.846016
Rwneg28_81 in28 sn81 11140.846016
Rwneg28_82 in28 sn82 11140.846016
Rwneg28_83 in28 sn83 11140.846016
Rwneg28_84 in28 sn84 11140.846016
Rwneg28_85 in28 sn85 3183.098862
Rwneg28_86 in28 sn86 3183.098862
Rwneg28_87 in28 sn87 11140.846016
Rwneg28_88 in28 sn88 3183.098862
Rwneg28_89 in28 sn89 11140.846016
Rwneg28_90 in28 sn90 3183.098862
Rwneg28_91 in28 sn91 3183.098862
Rwneg28_92 in28 sn92 3183.098862
Rwneg28_93 in28 sn93 11140.846016
Rwneg28_94 in28 sn94 3183.098862
Rwneg28_95 in28 sn95 3183.098862
Rwneg28_96 in28 sn96 11140.846016
Rwneg28_97 in28 sn97 11140.846016
Rwneg28_98 in28 sn98 11140.846016
Rwneg28_99 in28 sn99 3183.098862
Rwneg28_100 in28 sn100 3183.098862
Rwneg29_1 in29 sn1 11140.846016
Rwneg29_2 in29 sn2 11140.846016
Rwneg29_3 in29 sn3 11140.846016
Rwneg29_4 in29 sn4 3183.098862
Rwneg29_5 in29 sn5 3183.098862
Rwneg29_6 in29 sn6 3183.098862
Rwneg29_7 in29 sn7 11140.846016
Rwneg29_8 in29 sn8 11140.846016
Rwneg29_9 in29 sn9 11140.846016
Rwneg29_10 in29 sn10 3183.098862
Rwneg29_11 in29 sn11 3183.098862
Rwneg29_12 in29 sn12 3183.098862
Rwneg29_13 in29 sn13 11140.846016
Rwneg29_14 in29 sn14 11140.846016
Rwneg29_15 in29 sn15 11140.846016
Rwneg29_16 in29 sn16 3183.098862
Rwneg29_17 in29 sn17 3183.098862
Rwneg29_18 in29 sn18 3183.098862
Rwneg29_19 in29 sn19 11140.846016
Rwneg29_20 in29 sn20 11140.846016
Rwneg29_21 in29 sn21 11140.846016
Rwneg29_22 in29 sn22 11140.846016
Rwneg29_23 in29 sn23 11140.846016
Rwneg29_24 in29 sn24 11140.846016
Rwneg29_25 in29 sn25 11140.846016
Rwneg29_26 in29 sn26 11140.846016
Rwneg29_27 in29 sn27 3183.098862
Rwneg29_28 in29 sn28 11140.846016
Rwneg29_29 in29 sn29 3183.098862
Rwneg29_30 in29 sn30 3183.098862
Rwneg29_31 in29 sn31 3183.098862
Rwneg29_32 in29 sn32 3183.098862
Rwneg29_33 in29 sn33 3183.098862
Rwneg29_34 in29 sn34 11140.846016
Rwneg29_35 in29 sn35 11140.846016
Rwneg29_36 in29 sn36 3183.098862
Rwneg29_37 in29 sn37 3183.098862
Rwneg29_38 in29 sn38 3183.098862
Rwneg29_39 in29 sn39 11140.846016
Rwneg29_40 in29 sn40 11140.846016
Rwneg29_41 in29 sn41 11140.846016
Rwneg29_42 in29 sn42 3183.098862
Rwneg29_43 in29 sn43 3183.098862
Rwneg29_44 in29 sn44 11140.846016
Rwneg29_45 in29 sn45 11140.846016
Rwneg29_46 in29 sn46 11140.846016
Rwneg29_47 in29 sn47 11140.846016
Rwneg29_48 in29 sn48 3183.098862
Rwneg29_49 in29 sn49 3183.098862
Rwneg29_50 in29 sn50 11140.846016
Rwneg29_51 in29 sn51 11140.846016
Rwneg29_52 in29 sn52 11140.846016
Rwneg29_53 in29 sn53 3183.098862
Rwneg29_54 in29 sn54 3183.098862
Rwneg29_55 in29 sn55 11140.846016
Rwneg29_56 in29 sn56 11140.846016
Rwneg29_57 in29 sn57 11140.846016
Rwneg29_58 in29 sn58 11140.846016
Rwneg29_59 in29 sn59 3183.098862
Rwneg29_60 in29 sn60 11140.846016
Rwneg29_61 in29 sn61 3183.098862
Rwneg29_62 in29 sn62 11140.846016
Rwneg29_63 in29 sn63 11140.846016
Rwneg29_64 in29 sn64 11140.846016
Rwneg29_65 in29 sn65 3183.098862
Rwneg29_66 in29 sn66 3183.098862
Rwneg29_67 in29 sn67 11140.846016
Rwneg29_68 in29 sn68 3183.098862
Rwneg29_69 in29 sn69 3183.098862
Rwneg29_70 in29 sn70 3183.098862
Rwneg29_71 in29 sn71 11140.846016
Rwneg29_72 in29 sn72 11140.846016
Rwneg29_73 in29 sn73 11140.846016
Rwneg29_74 in29 sn74 11140.846016
Rwneg29_75 in29 sn75 3183.098862
Rwneg29_76 in29 sn76 3183.098862
Rwneg29_77 in29 sn77 11140.846016
Rwneg29_78 in29 sn78 3183.098862
Rwneg29_79 in29 sn79 3183.098862
Rwneg29_80 in29 sn80 11140.846016
Rwneg29_81 in29 sn81 3183.098862
Rwneg29_82 in29 sn82 3183.098862
Rwneg29_83 in29 sn83 3183.098862
Rwneg29_84 in29 sn84 3183.098862
Rwneg29_85 in29 sn85 11140.846016
Rwneg29_86 in29 sn86 3183.098862
Rwneg29_87 in29 sn87 11140.846016
Rwneg29_88 in29 sn88 11140.846016
Rwneg29_89 in29 sn89 11140.846016
Rwneg29_90 in29 sn90 11140.846016
Rwneg29_91 in29 sn91 3183.098862
Rwneg29_92 in29 sn92 3183.098862
Rwneg29_93 in29 sn93 11140.846016
Rwneg29_94 in29 sn94 11140.846016
Rwneg29_95 in29 sn95 11140.846016
Rwneg29_96 in29 sn96 3183.098862
Rwneg29_97 in29 sn97 11140.846016
Rwneg29_98 in29 sn98 11140.846016
Rwneg29_99 in29 sn99 3183.098862
Rwneg29_100 in29 sn100 11140.846016
Rwneg30_1 in30 sn1 3183.098862
Rwneg30_2 in30 sn2 3183.098862
Rwneg30_3 in30 sn3 11140.846016
Rwneg30_4 in30 sn4 11140.846016
Rwneg30_5 in30 sn5 11140.846016
Rwneg30_6 in30 sn6 11140.846016
Rwneg30_7 in30 sn7 3183.098862
Rwneg30_8 in30 sn8 3183.098862
Rwneg30_9 in30 sn9 3183.098862
Rwneg30_10 in30 sn10 11140.846016
Rwneg30_11 in30 sn11 11140.846016
Rwneg30_12 in30 sn12 3183.098862
Rwneg30_13 in30 sn13 3183.098862
Rwneg30_14 in30 sn14 11140.846016
Rwneg30_15 in30 sn15 3183.098862
Rwneg30_16 in30 sn16 3183.098862
Rwneg30_17 in30 sn17 11140.846016
Rwneg30_18 in30 sn18 3183.098862
Rwneg30_19 in30 sn19 11140.846016
Rwneg30_20 in30 sn20 11140.846016
Rwneg30_21 in30 sn21 3183.098862
Rwneg30_22 in30 sn22 11140.846016
Rwneg30_23 in30 sn23 3183.098862
Rwneg30_24 in30 sn24 11140.846016
Rwneg30_25 in30 sn25 11140.846016
Rwneg30_26 in30 sn26 3183.098862
Rwneg30_27 in30 sn27 11140.846016
Rwneg30_28 in30 sn28 11140.846016
Rwneg30_29 in30 sn29 3183.098862
Rwneg30_30 in30 sn30 11140.846016
Rwneg30_31 in30 sn31 3183.098862
Rwneg30_32 in30 sn32 11140.846016
Rwneg30_33 in30 sn33 11140.846016
Rwneg30_34 in30 sn34 11140.846016
Rwneg30_35 in30 sn35 11140.846016
Rwneg30_36 in30 sn36 3183.098862
Rwneg30_37 in30 sn37 3183.098862
Rwneg30_38 in30 sn38 11140.846016
Rwneg30_39 in30 sn39 3183.098862
Rwneg30_40 in30 sn40 3183.098862
Rwneg30_41 in30 sn41 3183.098862
Rwneg30_42 in30 sn42 11140.846016
Rwneg30_43 in30 sn43 3183.098862
Rwneg30_44 in30 sn44 3183.098862
Rwneg30_45 in30 sn45 3183.098862
Rwneg30_46 in30 sn46 11140.846016
Rwneg30_47 in30 sn47 3183.098862
Rwneg30_48 in30 sn48 11140.846016
Rwneg30_49 in30 sn49 11140.846016
Rwneg30_50 in30 sn50 3183.098862
Rwneg30_51 in30 sn51 11140.846016
Rwneg30_52 in30 sn52 11140.846016
Rwneg30_53 in30 sn53 11140.846016
Rwneg30_54 in30 sn54 11140.846016
Rwneg30_55 in30 sn55 3183.098862
Rwneg30_56 in30 sn56 3183.098862
Rwneg30_57 in30 sn57 11140.846016
Rwneg30_58 in30 sn58 3183.098862
Rwneg30_59 in30 sn59 3183.098862
Rwneg30_60 in30 sn60 11140.846016
Rwneg30_61 in30 sn61 11140.846016
Rwneg30_62 in30 sn62 11140.846016
Rwneg30_63 in30 sn63 3183.098862
Rwneg30_64 in30 sn64 11140.846016
Rwneg30_65 in30 sn65 3183.098862
Rwneg30_66 in30 sn66 3183.098862
Rwneg30_67 in30 sn67 11140.846016
Rwneg30_68 in30 sn68 3183.098862
Rwneg30_69 in30 sn69 11140.846016
Rwneg30_70 in30 sn70 11140.846016
Rwneg30_71 in30 sn71 3183.098862
Rwneg30_72 in30 sn72 3183.098862
Rwneg30_73 in30 sn73 3183.098862
Rwneg30_74 in30 sn74 3183.098862
Rwneg30_75 in30 sn75 3183.098862
Rwneg30_76 in30 sn76 11140.846016
Rwneg30_77 in30 sn77 3183.098862
Rwneg30_78 in30 sn78 11140.846016
Rwneg30_79 in30 sn79 3183.098862
Rwneg30_80 in30 sn80 11140.846016
Rwneg30_81 in30 sn81 3183.098862
Rwneg30_82 in30 sn82 3183.098862
Rwneg30_83 in30 sn83 11140.846016
Rwneg30_84 in30 sn84 11140.846016
Rwneg30_85 in30 sn85 11140.846016
Rwneg30_86 in30 sn86 11140.846016
Rwneg30_87 in30 sn87 3183.098862
Rwneg30_88 in30 sn88 11140.846016
Rwneg30_89 in30 sn89 11140.846016
Rwneg30_90 in30 sn90 11140.846016
Rwneg30_91 in30 sn91 11140.846016
Rwneg30_92 in30 sn92 11140.846016
Rwneg30_93 in30 sn93 11140.846016
Rwneg30_94 in30 sn94 3183.098862
Rwneg30_95 in30 sn95 3183.098862
Rwneg30_96 in30 sn96 3183.098862
Rwneg30_97 in30 sn97 11140.846016
Rwneg30_98 in30 sn98 11140.846016
Rwneg30_99 in30 sn99 3183.098862
Rwneg30_100 in30 sn100 11140.846016
Rwneg31_1 in31 sn1 11140.846016
Rwneg31_2 in31 sn2 3183.098862
Rwneg31_3 in31 sn3 3183.098862
Rwneg31_4 in31 sn4 3183.098862
Rwneg31_5 in31 sn5 3183.098862
Rwneg31_6 in31 sn6 3183.098862
Rwneg31_7 in31 sn7 3183.098862
Rwneg31_8 in31 sn8 11140.846016
Rwneg31_9 in31 sn9 11140.846016
Rwneg31_10 in31 sn10 3183.098862
Rwneg31_11 in31 sn11 11140.846016
Rwneg31_12 in31 sn12 11140.846016
Rwneg31_13 in31 sn13 3183.098862
Rwneg31_14 in31 sn14 11140.846016
Rwneg31_15 in31 sn15 3183.098862
Rwneg31_16 in31 sn16 11140.846016
Rwneg31_17 in31 sn17 11140.846016
Rwneg31_18 in31 sn18 3183.098862
Rwneg31_19 in31 sn19 11140.846016
Rwneg31_20 in31 sn20 11140.846016
Rwneg31_21 in31 sn21 11140.846016
Rwneg31_22 in31 sn22 3183.098862
Rwneg31_23 in31 sn23 11140.846016
Rwneg31_24 in31 sn24 11140.846016
Rwneg31_25 in31 sn25 3183.098862
Rwneg31_26 in31 sn26 3183.098862
Rwneg31_27 in31 sn27 11140.846016
Rwneg31_28 in31 sn28 11140.846016
Rwneg31_29 in31 sn29 3183.098862
Rwneg31_30 in31 sn30 11140.846016
Rwneg31_31 in31 sn31 3183.098862
Rwneg31_32 in31 sn32 3183.098862
Rwneg31_33 in31 sn33 3183.098862
Rwneg31_34 in31 sn34 11140.846016
Rwneg31_35 in31 sn35 11140.846016
Rwneg31_36 in31 sn36 3183.098862
Rwneg31_37 in31 sn37 11140.846016
Rwneg31_38 in31 sn38 11140.846016
Rwneg31_39 in31 sn39 3183.098862
Rwneg31_40 in31 sn40 11140.846016
Rwneg31_41 in31 sn41 11140.846016
Rwneg31_42 in31 sn42 3183.098862
Rwneg31_43 in31 sn43 11140.846016
Rwneg31_44 in31 sn44 3183.098862
Rwneg31_45 in31 sn45 11140.846016
Rwneg31_46 in31 sn46 11140.846016
Rwneg31_47 in31 sn47 3183.098862
Rwneg31_48 in31 sn48 11140.846016
Rwneg31_49 in31 sn49 3183.098862
Rwneg31_50 in31 sn50 3183.098862
Rwneg31_51 in31 sn51 11140.846016
Rwneg31_52 in31 sn52 3183.098862
Rwneg31_53 in31 sn53 3183.098862
Rwneg31_54 in31 sn54 11140.846016
Rwneg31_55 in31 sn55 11140.846016
Rwneg31_56 in31 sn56 11140.846016
Rwneg31_57 in31 sn57 11140.846016
Rwneg31_58 in31 sn58 3183.098862
Rwneg31_59 in31 sn59 11140.846016
Rwneg31_60 in31 sn60 11140.846016
Rwneg31_61 in31 sn61 11140.846016
Rwneg31_62 in31 sn62 11140.846016
Rwneg31_63 in31 sn63 3183.098862
Rwneg31_64 in31 sn64 3183.098862
Rwneg31_65 in31 sn65 3183.098862
Rwneg31_66 in31 sn66 3183.098862
Rwneg31_67 in31 sn67 11140.846016
Rwneg31_68 in31 sn68 11140.846016
Rwneg31_69 in31 sn69 3183.098862
Rwneg31_70 in31 sn70 11140.846016
Rwneg31_71 in31 sn71 3183.098862
Rwneg31_72 in31 sn72 11140.846016
Rwneg31_73 in31 sn73 11140.846016
Rwneg31_74 in31 sn74 11140.846016
Rwneg31_75 in31 sn75 11140.846016
Rwneg31_76 in31 sn76 11140.846016
Rwneg31_77 in31 sn77 11140.846016
Rwneg31_78 in31 sn78 11140.846016
Rwneg31_79 in31 sn79 3183.098862
Rwneg31_80 in31 sn80 11140.846016
Rwneg31_81 in31 sn81 3183.098862
Rwneg31_82 in31 sn82 11140.846016
Rwneg31_83 in31 sn83 3183.098862
Rwneg31_84 in31 sn84 11140.846016
Rwneg31_85 in31 sn85 3183.098862
Rwneg31_86 in31 sn86 11140.846016
Rwneg31_87 in31 sn87 11140.846016
Rwneg31_88 in31 sn88 11140.846016
Rwneg31_89 in31 sn89 3183.098862
Rwneg31_90 in31 sn90 11140.846016
Rwneg31_91 in31 sn91 11140.846016
Rwneg31_92 in31 sn92 11140.846016
Rwneg31_93 in31 sn93 3183.098862
Rwneg31_94 in31 sn94 3183.098862
Rwneg31_95 in31 sn95 3183.098862
Rwneg31_96 in31 sn96 3183.098862
Rwneg31_97 in31 sn97 11140.846016
Rwneg31_98 in31 sn98 11140.846016
Rwneg31_99 in31 sn99 3183.098862
Rwneg31_100 in31 sn100 11140.846016
Rwneg32_1 in32 sn1 3183.098862
Rwneg32_2 in32 sn2 11140.846016
Rwneg32_3 in32 sn3 11140.846016
Rwneg32_4 in32 sn4 3183.098862
Rwneg32_5 in32 sn5 3183.098862
Rwneg32_6 in32 sn6 3183.098862
Rwneg32_7 in32 sn7 11140.846016
Rwneg32_8 in32 sn8 11140.846016
Rwneg32_9 in32 sn9 11140.846016
Rwneg32_10 in32 sn10 11140.846016
Rwneg32_11 in32 sn11 3183.098862
Rwneg32_12 in32 sn12 3183.098862
Rwneg32_13 in32 sn13 11140.846016
Rwneg32_14 in32 sn14 11140.846016
Rwneg32_15 in32 sn15 3183.098862
Rwneg32_16 in32 sn16 11140.846016
Rwneg32_17 in32 sn17 3183.098862
Rwneg32_18 in32 sn18 11140.846016
Rwneg32_19 in32 sn19 11140.846016
Rwneg32_20 in32 sn20 3183.098862
Rwneg32_21 in32 sn21 11140.846016
Rwneg32_22 in32 sn22 11140.846016
Rwneg32_23 in32 sn23 11140.846016
Rwneg32_24 in32 sn24 3183.098862
Rwneg32_25 in32 sn25 3183.098862
Rwneg32_26 in32 sn26 3183.098862
Rwneg32_27 in32 sn27 3183.098862
Rwneg32_28 in32 sn28 11140.846016
Rwneg32_29 in32 sn29 11140.846016
Rwneg32_30 in32 sn30 11140.846016
Rwneg32_31 in32 sn31 11140.846016
Rwneg32_32 in32 sn32 3183.098862
Rwneg32_33 in32 sn33 11140.846016
Rwneg32_34 in32 sn34 3183.098862
Rwneg32_35 in32 sn35 3183.098862
Rwneg32_36 in32 sn36 11140.846016
Rwneg32_37 in32 sn37 11140.846016
Rwneg32_38 in32 sn38 3183.098862
Rwneg32_39 in32 sn39 11140.846016
Rwneg32_40 in32 sn40 11140.846016
Rwneg32_41 in32 sn41 11140.846016
Rwneg32_42 in32 sn42 11140.846016
Rwneg32_43 in32 sn43 11140.846016
Rwneg32_44 in32 sn44 11140.846016
Rwneg32_45 in32 sn45 3183.098862
Rwneg32_46 in32 sn46 3183.098862
Rwneg32_47 in32 sn47 11140.846016
Rwneg32_48 in32 sn48 11140.846016
Rwneg32_49 in32 sn49 3183.098862
Rwneg32_50 in32 sn50 3183.098862
Rwneg32_51 in32 sn51 3183.098862
Rwneg32_52 in32 sn52 3183.098862
Rwneg32_53 in32 sn53 11140.846016
Rwneg32_54 in32 sn54 11140.846016
Rwneg32_55 in32 sn55 11140.846016
Rwneg32_56 in32 sn56 11140.846016
Rwneg32_57 in32 sn57 3183.098862
Rwneg32_58 in32 sn58 3183.098862
Rwneg32_59 in32 sn59 11140.846016
Rwneg32_60 in32 sn60 3183.098862
Rwneg32_61 in32 sn61 3183.098862
Rwneg32_62 in32 sn62 11140.846016
Rwneg32_63 in32 sn63 3183.098862
Rwneg32_64 in32 sn64 11140.846016
Rwneg32_65 in32 sn65 3183.098862
Rwneg32_66 in32 sn66 11140.846016
Rwneg32_67 in32 sn67 11140.846016
Rwneg32_68 in32 sn68 11140.846016
Rwneg32_69 in32 sn69 11140.846016
Rwneg32_70 in32 sn70 3183.098862
Rwneg32_71 in32 sn71 3183.098862
Rwneg32_72 in32 sn72 3183.098862
Rwneg32_73 in32 sn73 3183.098862
Rwneg32_74 in32 sn74 11140.846016
Rwneg32_75 in32 sn75 11140.846016
Rwneg32_76 in32 sn76 3183.098862
Rwneg32_77 in32 sn77 11140.846016
Rwneg32_78 in32 sn78 3183.098862
Rwneg32_79 in32 sn79 3183.098862
Rwneg32_80 in32 sn80 11140.846016
Rwneg32_81 in32 sn81 3183.098862
Rwneg32_82 in32 sn82 11140.846016
Rwneg32_83 in32 sn83 11140.846016
Rwneg32_84 in32 sn84 11140.846016
Rwneg32_85 in32 sn85 3183.098862
Rwneg32_86 in32 sn86 3183.098862
Rwneg32_87 in32 sn87 11140.846016
Rwneg32_88 in32 sn88 11140.846016
Rwneg32_89 in32 sn89 3183.098862
Rwneg32_90 in32 sn90 3183.098862
Rwneg32_91 in32 sn91 11140.846016
Rwneg32_92 in32 sn92 3183.098862
Rwneg32_93 in32 sn93 11140.846016
Rwneg32_94 in32 sn94 11140.846016
Rwneg32_95 in32 sn95 3183.098862
Rwneg32_96 in32 sn96 3183.098862
Rwneg32_97 in32 sn97 3183.098862
Rwneg32_98 in32 sn98 11140.846016
Rwneg32_99 in32 sn99 11140.846016
Rwneg32_100 in32 sn100 3183.098862
Rwneg33_1 in33 sn1 3183.098862
Rwneg33_2 in33 sn2 11140.846016
Rwneg33_3 in33 sn3 3183.098862
Rwneg33_4 in33 sn4 3183.098862
Rwneg33_5 in33 sn5 11140.846016
Rwneg33_6 in33 sn6 3183.098862
Rwneg33_7 in33 sn7 11140.846016
Rwneg33_8 in33 sn8 11140.846016
Rwneg33_9 in33 sn9 11140.846016
Rwneg33_10 in33 sn10 11140.846016
Rwneg33_11 in33 sn11 3183.098862
Rwneg33_12 in33 sn12 11140.846016
Rwneg33_13 in33 sn13 3183.098862
Rwneg33_14 in33 sn14 11140.846016
Rwneg33_15 in33 sn15 3183.098862
Rwneg33_16 in33 sn16 11140.846016
Rwneg33_17 in33 sn17 3183.098862
Rwneg33_18 in33 sn18 3183.098862
Rwneg33_19 in33 sn19 11140.846016
Rwneg33_20 in33 sn20 3183.098862
Rwneg33_21 in33 sn21 3183.098862
Rwneg33_22 in33 sn22 11140.846016
Rwneg33_23 in33 sn23 11140.846016
Rwneg33_24 in33 sn24 11140.846016
Rwneg33_25 in33 sn25 11140.846016
Rwneg33_26 in33 sn26 3183.098862
Rwneg33_27 in33 sn27 3183.098862
Rwneg33_28 in33 sn28 11140.846016
Rwneg33_29 in33 sn29 3183.098862
Rwneg33_30 in33 sn30 11140.846016
Rwneg33_31 in33 sn31 3183.098862
Rwneg33_32 in33 sn32 11140.846016
Rwneg33_33 in33 sn33 3183.098862
Rwneg33_34 in33 sn34 3183.098862
Rwneg33_35 in33 sn35 11140.846016
Rwneg33_36 in33 sn36 3183.098862
Rwneg33_37 in33 sn37 3183.098862
Rwneg33_38 in33 sn38 3183.098862
Rwneg33_39 in33 sn39 3183.098862
Rwneg33_40 in33 sn40 11140.846016
Rwneg33_41 in33 sn41 3183.098862
Rwneg33_42 in33 sn42 3183.098862
Rwneg33_43 in33 sn43 3183.098862
Rwneg33_44 in33 sn44 3183.098862
Rwneg33_45 in33 sn45 3183.098862
Rwneg33_46 in33 sn46 3183.098862
Rwneg33_47 in33 sn47 3183.098862
Rwneg33_48 in33 sn48 11140.846016
Rwneg33_49 in33 sn49 3183.098862
Rwneg33_50 in33 sn50 11140.846016
Rwneg33_51 in33 sn51 11140.846016
Rwneg33_52 in33 sn52 3183.098862
Rwneg33_53 in33 sn53 3183.098862
Rwneg33_54 in33 sn54 3183.098862
Rwneg33_55 in33 sn55 11140.846016
Rwneg33_56 in33 sn56 3183.098862
Rwneg33_57 in33 sn57 11140.846016
Rwneg33_58 in33 sn58 3183.098862
Rwneg33_59 in33 sn59 3183.098862
Rwneg33_60 in33 sn60 11140.846016
Rwneg33_61 in33 sn61 11140.846016
Rwneg33_62 in33 sn62 11140.846016
Rwneg33_63 in33 sn63 3183.098862
Rwneg33_64 in33 sn64 11140.846016
Rwneg33_65 in33 sn65 3183.098862
Rwneg33_66 in33 sn66 3183.098862
Rwneg33_67 in33 sn67 11140.846016
Rwneg33_68 in33 sn68 3183.098862
Rwneg33_69 in33 sn69 11140.846016
Rwneg33_70 in33 sn70 11140.846016
Rwneg33_71 in33 sn71 11140.846016
Rwneg33_72 in33 sn72 11140.846016
Rwneg33_73 in33 sn73 11140.846016
Rwneg33_74 in33 sn74 11140.846016
Rwneg33_75 in33 sn75 3183.098862
Rwneg33_76 in33 sn76 3183.098862
Rwneg33_77 in33 sn77 11140.846016
Rwneg33_78 in33 sn78 11140.846016
Rwneg33_79 in33 sn79 11140.846016
Rwneg33_80 in33 sn80 3183.098862
Rwneg33_81 in33 sn81 3183.098862
Rwneg33_82 in33 sn82 3183.098862
Rwneg33_83 in33 sn83 11140.846016
Rwneg33_84 in33 sn84 11140.846016
Rwneg33_85 in33 sn85 3183.098862
Rwneg33_86 in33 sn86 3183.098862
Rwneg33_87 in33 sn87 11140.846016
Rwneg33_88 in33 sn88 3183.098862
Rwneg33_89 in33 sn89 3183.098862
Rwneg33_90 in33 sn90 11140.846016
Rwneg33_91 in33 sn91 3183.098862
Rwneg33_92 in33 sn92 11140.846016
Rwneg33_93 in33 sn93 11140.846016
Rwneg33_94 in33 sn94 11140.846016
Rwneg33_95 in33 sn95 3183.098862
Rwneg33_96 in33 sn96 11140.846016
Rwneg33_97 in33 sn97 3183.098862
Rwneg33_98 in33 sn98 3183.098862
Rwneg33_99 in33 sn99 11140.846016
Rwneg33_100 in33 sn100 3183.098862
Rwneg34_1 in34 sn1 11140.846016
Rwneg34_2 in34 sn2 11140.846016
Rwneg34_3 in34 sn3 11140.846016
Rwneg34_4 in34 sn4 11140.846016
Rwneg34_5 in34 sn5 3183.098862
Rwneg34_6 in34 sn6 3183.098862
Rwneg34_7 in34 sn7 3183.098862
Rwneg34_8 in34 sn8 3183.098862
Rwneg34_9 in34 sn9 3183.098862
Rwneg34_10 in34 sn10 3183.098862
Rwneg34_11 in34 sn11 3183.098862
Rwneg34_12 in34 sn12 3183.098862
Rwneg34_13 in34 sn13 11140.846016
Rwneg34_14 in34 sn14 11140.846016
Rwneg34_15 in34 sn15 3183.098862
Rwneg34_16 in34 sn16 3183.098862
Rwneg34_17 in34 sn17 11140.846016
Rwneg34_18 in34 sn18 11140.846016
Rwneg34_19 in34 sn19 11140.846016
Rwneg34_20 in34 sn20 11140.846016
Rwneg34_21 in34 sn21 3183.098862
Rwneg34_22 in34 sn22 11140.846016
Rwneg34_23 in34 sn23 3183.098862
Rwneg34_24 in34 sn24 11140.846016
Rwneg34_25 in34 sn25 3183.098862
Rwneg34_26 in34 sn26 11140.846016
Rwneg34_27 in34 sn27 3183.098862
Rwneg34_28 in34 sn28 3183.098862
Rwneg34_29 in34 sn29 3183.098862
Rwneg34_30 in34 sn30 11140.846016
Rwneg34_31 in34 sn31 3183.098862
Rwneg34_32 in34 sn32 11140.846016
Rwneg34_33 in34 sn33 11140.846016
Rwneg34_34 in34 sn34 11140.846016
Rwneg34_35 in34 sn35 3183.098862
Rwneg34_36 in34 sn36 3183.098862
Rwneg34_37 in34 sn37 3183.098862
Rwneg34_38 in34 sn38 11140.846016
Rwneg34_39 in34 sn39 11140.846016
Rwneg34_40 in34 sn40 3183.098862
Rwneg34_41 in34 sn41 11140.846016
Rwneg34_42 in34 sn42 3183.098862
Rwneg34_43 in34 sn43 3183.098862
Rwneg34_44 in34 sn44 11140.846016
Rwneg34_45 in34 sn45 3183.098862
Rwneg34_46 in34 sn46 11140.846016
Rwneg34_47 in34 sn47 3183.098862
Rwneg34_48 in34 sn48 11140.846016
Rwneg34_49 in34 sn49 11140.846016
Rwneg34_50 in34 sn50 11140.846016
Rwneg34_51 in34 sn51 11140.846016
Rwneg34_52 in34 sn52 3183.098862
Rwneg34_53 in34 sn53 11140.846016
Rwneg34_54 in34 sn54 11140.846016
Rwneg34_55 in34 sn55 3183.098862
Rwneg34_56 in34 sn56 3183.098862
Rwneg34_57 in34 sn57 11140.846016
Rwneg34_58 in34 sn58 3183.098862
Rwneg34_59 in34 sn59 3183.098862
Rwneg34_60 in34 sn60 11140.846016
Rwneg34_61 in34 sn61 11140.846016
Rwneg34_62 in34 sn62 11140.846016
Rwneg34_63 in34 sn63 3183.098862
Rwneg34_64 in34 sn64 11140.846016
Rwneg34_65 in34 sn65 11140.846016
Rwneg34_66 in34 sn66 3183.098862
Rwneg34_67 in34 sn67 3183.098862
Rwneg34_68 in34 sn68 3183.098862
Rwneg34_69 in34 sn69 11140.846016
Rwneg34_70 in34 sn70 11140.846016
Rwneg34_71 in34 sn71 3183.098862
Rwneg34_72 in34 sn72 3183.098862
Rwneg34_73 in34 sn73 3183.098862
Rwneg34_74 in34 sn74 11140.846016
Rwneg34_75 in34 sn75 11140.846016
Rwneg34_76 in34 sn76 3183.098862
Rwneg34_77 in34 sn77 11140.846016
Rwneg34_78 in34 sn78 11140.846016
Rwneg34_79 in34 sn79 3183.098862
Rwneg34_80 in34 sn80 11140.846016
Rwneg34_81 in34 sn81 11140.846016
Rwneg34_82 in34 sn82 11140.846016
Rwneg34_83 in34 sn83 11140.846016
Rwneg34_84 in34 sn84 11140.846016
Rwneg34_85 in34 sn85 3183.098862
Rwneg34_86 in34 sn86 11140.846016
Rwneg34_87 in34 sn87 3183.098862
Rwneg34_88 in34 sn88 3183.098862
Rwneg34_89 in34 sn89 11140.846016
Rwneg34_90 in34 sn90 3183.098862
Rwneg34_91 in34 sn91 11140.846016
Rwneg34_92 in34 sn92 11140.846016
Rwneg34_93 in34 sn93 11140.846016
Rwneg34_94 in34 sn94 11140.846016
Rwneg34_95 in34 sn95 3183.098862
Rwneg34_96 in34 sn96 11140.846016
Rwneg34_97 in34 sn97 11140.846016
Rwneg34_98 in34 sn98 3183.098862
Rwneg34_99 in34 sn99 11140.846016
Rwneg34_100 in34 sn100 3183.098862
Rwneg35_1 in35 sn1 3183.098862
Rwneg35_2 in35 sn2 11140.846016
Rwneg35_3 in35 sn3 11140.846016
Rwneg35_4 in35 sn4 11140.846016
Rwneg35_5 in35 sn5 3183.098862
Rwneg35_6 in35 sn6 3183.098862
Rwneg35_7 in35 sn7 11140.846016
Rwneg35_8 in35 sn8 3183.098862
Rwneg35_9 in35 sn9 3183.098862
Rwneg35_10 in35 sn10 11140.846016
Rwneg35_11 in35 sn11 3183.098862
Rwneg35_12 in35 sn12 3183.098862
Rwneg35_13 in35 sn13 3183.098862
Rwneg35_14 in35 sn14 11140.846016
Rwneg35_15 in35 sn15 3183.098862
Rwneg35_16 in35 sn16 11140.846016
Rwneg35_17 in35 sn17 3183.098862
Rwneg35_18 in35 sn18 11140.846016
Rwneg35_19 in35 sn19 3183.098862
Rwneg35_20 in35 sn20 3183.098862
Rwneg35_21 in35 sn21 11140.846016
Rwneg35_22 in35 sn22 11140.846016
Rwneg35_23 in35 sn23 3183.098862
Rwneg35_24 in35 sn24 11140.846016
Rwneg35_25 in35 sn25 11140.846016
Rwneg35_26 in35 sn26 11140.846016
Rwneg35_27 in35 sn27 3183.098862
Rwneg35_28 in35 sn28 11140.846016
Rwneg35_29 in35 sn29 11140.846016
Rwneg35_30 in35 sn30 11140.846016
Rwneg35_31 in35 sn31 11140.846016
Rwneg35_32 in35 sn32 11140.846016
Rwneg35_33 in35 sn33 3183.098862
Rwneg35_34 in35 sn34 11140.846016
Rwneg35_35 in35 sn35 11140.846016
Rwneg35_36 in35 sn36 3183.098862
Rwneg35_37 in35 sn37 3183.098862
Rwneg35_38 in35 sn38 3183.098862
Rwneg35_39 in35 sn39 3183.098862
Rwneg35_40 in35 sn40 11140.846016
Rwneg35_41 in35 sn41 11140.846016
Rwneg35_42 in35 sn42 11140.846016
Rwneg35_43 in35 sn43 11140.846016
Rwneg35_44 in35 sn44 3183.098862
Rwneg35_45 in35 sn45 3183.098862
Rwneg35_46 in35 sn46 11140.846016
Rwneg35_47 in35 sn47 3183.098862
Rwneg35_48 in35 sn48 3183.098862
Rwneg35_49 in35 sn49 3183.098862
Rwneg35_50 in35 sn50 11140.846016
Rwneg35_51 in35 sn51 11140.846016
Rwneg35_52 in35 sn52 3183.098862
Rwneg35_53 in35 sn53 11140.846016
Rwneg35_54 in35 sn54 11140.846016
Rwneg35_55 in35 sn55 11140.846016
Rwneg35_56 in35 sn56 11140.846016
Rwneg35_57 in35 sn57 3183.098862
Rwneg35_58 in35 sn58 3183.098862
Rwneg35_59 in35 sn59 3183.098862
Rwneg35_60 in35 sn60 3183.098862
Rwneg35_61 in35 sn61 3183.098862
Rwneg35_62 in35 sn62 11140.846016
Rwneg35_63 in35 sn63 3183.098862
Rwneg35_64 in35 sn64 3183.098862
Rwneg35_65 in35 sn65 11140.846016
Rwneg35_66 in35 sn66 11140.846016
Rwneg35_67 in35 sn67 3183.098862
Rwneg35_68 in35 sn68 3183.098862
Rwneg35_69 in35 sn69 3183.098862
Rwneg35_70 in35 sn70 3183.098862
Rwneg35_71 in35 sn71 3183.098862
Rwneg35_72 in35 sn72 11140.846016
Rwneg35_73 in35 sn73 11140.846016
Rwneg35_74 in35 sn74 3183.098862
Rwneg35_75 in35 sn75 11140.846016
Rwneg35_76 in35 sn76 3183.098862
Rwneg35_77 in35 sn77 11140.846016
Rwneg35_78 in35 sn78 11140.846016
Rwneg35_79 in35 sn79 3183.098862
Rwneg35_80 in35 sn80 11140.846016
Rwneg35_81 in35 sn81 3183.098862
Rwneg35_82 in35 sn82 3183.098862
Rwneg35_83 in35 sn83 11140.846016
Rwneg35_84 in35 sn84 3183.098862
Rwneg35_85 in35 sn85 3183.098862
Rwneg35_86 in35 sn86 3183.098862
Rwneg35_87 in35 sn87 11140.846016
Rwneg35_88 in35 sn88 11140.846016
Rwneg35_89 in35 sn89 11140.846016
Rwneg35_90 in35 sn90 3183.098862
Rwneg35_91 in35 sn91 11140.846016
Rwneg35_92 in35 sn92 11140.846016
Rwneg35_93 in35 sn93 11140.846016
Rwneg35_94 in35 sn94 11140.846016
Rwneg35_95 in35 sn95 11140.846016
Rwneg35_96 in35 sn96 3183.098862
Rwneg35_97 in35 sn97 11140.846016
Rwneg35_98 in35 sn98 3183.098862
Rwneg35_99 in35 sn99 3183.098862
Rwneg35_100 in35 sn100 11140.846016
Rwneg36_1 in36 sn1 3183.098862
Rwneg36_2 in36 sn2 3183.098862
Rwneg36_3 in36 sn3 3183.098862
Rwneg36_4 in36 sn4 11140.846016
Rwneg36_5 in36 sn5 11140.846016
Rwneg36_6 in36 sn6 3183.098862
Rwneg36_7 in36 sn7 11140.846016
Rwneg36_8 in36 sn8 11140.846016
Rwneg36_9 in36 sn9 11140.846016
Rwneg36_10 in36 sn10 11140.846016
Rwneg36_11 in36 sn11 3183.098862
Rwneg36_12 in36 sn12 11140.846016
Rwneg36_13 in36 sn13 3183.098862
Rwneg36_14 in36 sn14 3183.098862
Rwneg36_15 in36 sn15 11140.846016
Rwneg36_16 in36 sn16 11140.846016
Rwneg36_17 in36 sn17 3183.098862
Rwneg36_18 in36 sn18 3183.098862
Rwneg36_19 in36 sn19 11140.846016
Rwneg36_20 in36 sn20 11140.846016
Rwneg36_21 in36 sn21 11140.846016
Rwneg36_22 in36 sn22 11140.846016
Rwneg36_23 in36 sn23 11140.846016
Rwneg36_24 in36 sn24 11140.846016
Rwneg36_25 in36 sn25 11140.846016
Rwneg36_26 in36 sn26 11140.846016
Rwneg36_27 in36 sn27 3183.098862
Rwneg36_28 in36 sn28 11140.846016
Rwneg36_29 in36 sn29 3183.098862
Rwneg36_30 in36 sn30 3183.098862
Rwneg36_31 in36 sn31 11140.846016
Rwneg36_32 in36 sn32 11140.846016
Rwneg36_33 in36 sn33 3183.098862
Rwneg36_34 in36 sn34 11140.846016
Rwneg36_35 in36 sn35 11140.846016
Rwneg36_36 in36 sn36 11140.846016
Rwneg36_37 in36 sn37 11140.846016
Rwneg36_38 in36 sn38 3183.098862
Rwneg36_39 in36 sn39 3183.098862
Rwneg36_40 in36 sn40 11140.846016
Rwneg36_41 in36 sn41 3183.098862
Rwneg36_42 in36 sn42 3183.098862
Rwneg36_43 in36 sn43 3183.098862
Rwneg36_44 in36 sn44 11140.846016
Rwneg36_45 in36 sn45 11140.846016
Rwneg36_46 in36 sn46 11140.846016
Rwneg36_47 in36 sn47 3183.098862
Rwneg36_48 in36 sn48 3183.098862
Rwneg36_49 in36 sn49 3183.098862
Rwneg36_50 in36 sn50 3183.098862
Rwneg36_51 in36 sn51 11140.846016
Rwneg36_52 in36 sn52 3183.098862
Rwneg36_53 in36 sn53 11140.846016
Rwneg36_54 in36 sn54 11140.846016
Rwneg36_55 in36 sn55 3183.098862
Rwneg36_56 in36 sn56 11140.846016
Rwneg36_57 in36 sn57 11140.846016
Rwneg36_58 in36 sn58 11140.846016
Rwneg36_59 in36 sn59 11140.846016
Rwneg36_60 in36 sn60 11140.846016
Rwneg36_61 in36 sn61 3183.098862
Rwneg36_62 in36 sn62 11140.846016
Rwneg36_63 in36 sn63 11140.846016
Rwneg36_64 in36 sn64 11140.846016
Rwneg36_65 in36 sn65 3183.098862
Rwneg36_66 in36 sn66 11140.846016
Rwneg36_67 in36 sn67 3183.098862
Rwneg36_68 in36 sn68 11140.846016
Rwneg36_69 in36 sn69 3183.098862
Rwneg36_70 in36 sn70 3183.098862
Rwneg36_71 in36 sn71 11140.846016
Rwneg36_72 in36 sn72 11140.846016
Rwneg36_73 in36 sn73 11140.846016
Rwneg36_74 in36 sn74 3183.098862
Rwneg36_75 in36 sn75 11140.846016
Rwneg36_76 in36 sn76 3183.098862
Rwneg36_77 in36 sn77 11140.846016
Rwneg36_78 in36 sn78 11140.846016
Rwneg36_79 in36 sn79 11140.846016
Rwneg36_80 in36 sn80 11140.846016
Rwneg36_81 in36 sn81 3183.098862
Rwneg36_82 in36 sn82 11140.846016
Rwneg36_83 in36 sn83 11140.846016
Rwneg36_84 in36 sn84 11140.846016
Rwneg36_85 in36 sn85 11140.846016
Rwneg36_86 in36 sn86 11140.846016
Rwneg36_87 in36 sn87 3183.098862
Rwneg36_88 in36 sn88 3183.098862
Rwneg36_89 in36 sn89 3183.098862
Rwneg36_90 in36 sn90 3183.098862
Rwneg36_91 in36 sn91 11140.846016
Rwneg36_92 in36 sn92 11140.846016
Rwneg36_93 in36 sn93 11140.846016
Rwneg36_94 in36 sn94 11140.846016
Rwneg36_95 in36 sn95 3183.098862
Rwneg36_96 in36 sn96 11140.846016
Rwneg36_97 in36 sn97 11140.846016
Rwneg36_98 in36 sn98 3183.098862
Rwneg36_99 in36 sn99 3183.098862
Rwneg36_100 in36 sn100 3183.098862
Rwneg37_1 in37 sn1 11140.846016
Rwneg37_2 in37 sn2 11140.846016
Rwneg37_3 in37 sn3 3183.098862
Rwneg37_4 in37 sn4 3183.098862
Rwneg37_5 in37 sn5 11140.846016
Rwneg37_6 in37 sn6 3183.098862
Rwneg37_7 in37 sn7 11140.846016
Rwneg37_8 in37 sn8 11140.846016
Rwneg37_9 in37 sn9 11140.846016
Rwneg37_10 in37 sn10 3183.098862
Rwneg37_11 in37 sn11 11140.846016
Rwneg37_12 in37 sn12 3183.098862
Rwneg37_13 in37 sn13 3183.098862
Rwneg37_14 in37 sn14 11140.846016
Rwneg37_15 in37 sn15 11140.846016
Rwneg37_16 in37 sn16 3183.098862
Rwneg37_17 in37 sn17 11140.846016
Rwneg37_18 in37 sn18 3183.098862
Rwneg37_19 in37 sn19 3183.098862
Rwneg37_20 in37 sn20 11140.846016
Rwneg37_21 in37 sn21 3183.098862
Rwneg37_22 in37 sn22 11140.846016
Rwneg37_23 in37 sn23 3183.098862
Rwneg37_24 in37 sn24 3183.098862
Rwneg37_25 in37 sn25 3183.098862
Rwneg37_26 in37 sn26 11140.846016
Rwneg37_27 in37 sn27 3183.098862
Rwneg37_28 in37 sn28 3183.098862
Rwneg37_29 in37 sn29 11140.846016
Rwneg37_30 in37 sn30 3183.098862
Rwneg37_31 in37 sn31 3183.098862
Rwneg37_32 in37 sn32 3183.098862
Rwneg37_33 in37 sn33 3183.098862
Rwneg37_34 in37 sn34 11140.846016
Rwneg37_35 in37 sn35 3183.098862
Rwneg37_36 in37 sn36 11140.846016
Rwneg37_37 in37 sn37 3183.098862
Rwneg37_38 in37 sn38 3183.098862
Rwneg37_39 in37 sn39 3183.098862
Rwneg37_40 in37 sn40 11140.846016
Rwneg37_41 in37 sn41 11140.846016
Rwneg37_42 in37 sn42 3183.098862
Rwneg37_43 in37 sn43 3183.098862
Rwneg37_44 in37 sn44 3183.098862
Rwneg37_45 in37 sn45 3183.098862
Rwneg37_46 in37 sn46 11140.846016
Rwneg37_47 in37 sn47 11140.846016
Rwneg37_48 in37 sn48 11140.846016
Rwneg37_49 in37 sn49 11140.846016
Rwneg37_50 in37 sn50 3183.098862
Rwneg37_51 in37 sn51 11140.846016
Rwneg37_52 in37 sn52 11140.846016
Rwneg37_53 in37 sn53 11140.846016
Rwneg37_54 in37 sn54 3183.098862
Rwneg37_55 in37 sn55 3183.098862
Rwneg37_56 in37 sn56 3183.098862
Rwneg37_57 in37 sn57 11140.846016
Rwneg37_58 in37 sn58 11140.846016
Rwneg37_59 in37 sn59 11140.846016
Rwneg37_60 in37 sn60 11140.846016
Rwneg37_61 in37 sn61 3183.098862
Rwneg37_62 in37 sn62 11140.846016
Rwneg37_63 in37 sn63 3183.098862
Rwneg37_64 in37 sn64 11140.846016
Rwneg37_65 in37 sn65 3183.098862
Rwneg37_66 in37 sn66 3183.098862
Rwneg37_67 in37 sn67 11140.846016
Rwneg37_68 in37 sn68 11140.846016
Rwneg37_69 in37 sn69 11140.846016
Rwneg37_70 in37 sn70 11140.846016
Rwneg37_71 in37 sn71 11140.846016
Rwneg37_72 in37 sn72 3183.098862
Rwneg37_73 in37 sn73 11140.846016
Rwneg37_74 in37 sn74 11140.846016
Rwneg37_75 in37 sn75 3183.098862
Rwneg37_76 in37 sn76 11140.846016
Rwneg37_77 in37 sn77 11140.846016
Rwneg37_78 in37 sn78 3183.098862
Rwneg37_79 in37 sn79 3183.098862
Rwneg37_80 in37 sn80 3183.098862
Rwneg37_81 in37 sn81 3183.098862
Rwneg37_82 in37 sn82 11140.846016
Rwneg37_83 in37 sn83 11140.846016
Rwneg37_84 in37 sn84 3183.098862
Rwneg37_85 in37 sn85 3183.098862
Rwneg37_86 in37 sn86 11140.846016
Rwneg37_87 in37 sn87 11140.846016
Rwneg37_88 in37 sn88 11140.846016
Rwneg37_89 in37 sn89 3183.098862
Rwneg37_90 in37 sn90 11140.846016
Rwneg37_91 in37 sn91 3183.098862
Rwneg37_92 in37 sn92 11140.846016
Rwneg37_93 in37 sn93 11140.846016
Rwneg37_94 in37 sn94 11140.846016
Rwneg37_95 in37 sn95 11140.846016
Rwneg37_96 in37 sn96 11140.846016
Rwneg37_97 in37 sn97 3183.098862
Rwneg37_98 in37 sn98 3183.098862
Rwneg37_99 in37 sn99 11140.846016
Rwneg37_100 in37 sn100 3183.098862
Rwneg38_1 in38 sn1 3183.098862
Rwneg38_2 in38 sn2 11140.846016
Rwneg38_3 in38 sn3 11140.846016
Rwneg38_4 in38 sn4 11140.846016
Rwneg38_5 in38 sn5 11140.846016
Rwneg38_6 in38 sn6 3183.098862
Rwneg38_7 in38 sn7 3183.098862
Rwneg38_8 in38 sn8 3183.098862
Rwneg38_9 in38 sn9 3183.098862
Rwneg38_10 in38 sn10 11140.846016
Rwneg38_11 in38 sn11 11140.846016
Rwneg38_12 in38 sn12 11140.846016
Rwneg38_13 in38 sn13 11140.846016
Rwneg38_14 in38 sn14 11140.846016
Rwneg38_15 in38 sn15 11140.846016
Rwneg38_16 in38 sn16 3183.098862
Rwneg38_17 in38 sn17 3183.098862
Rwneg38_18 in38 sn18 11140.846016
Rwneg38_19 in38 sn19 11140.846016
Rwneg38_20 in38 sn20 3183.098862
Rwneg38_21 in38 sn21 11140.846016
Rwneg38_22 in38 sn22 3183.098862
Rwneg38_23 in38 sn23 11140.846016
Rwneg38_24 in38 sn24 3183.098862
Rwneg38_25 in38 sn25 3183.098862
Rwneg38_26 in38 sn26 3183.098862
Rwneg38_27 in38 sn27 3183.098862
Rwneg38_28 in38 sn28 3183.098862
Rwneg38_29 in38 sn29 11140.846016
Rwneg38_30 in38 sn30 3183.098862
Rwneg38_31 in38 sn31 11140.846016
Rwneg38_32 in38 sn32 3183.098862
Rwneg38_33 in38 sn33 3183.098862
Rwneg38_34 in38 sn34 11140.846016
Rwneg38_35 in38 sn35 11140.846016
Rwneg38_36 in38 sn36 11140.846016
Rwneg38_37 in38 sn37 11140.846016
Rwneg38_38 in38 sn38 11140.846016
Rwneg38_39 in38 sn39 11140.846016
Rwneg38_40 in38 sn40 11140.846016
Rwneg38_41 in38 sn41 3183.098862
Rwneg38_42 in38 sn42 11140.846016
Rwneg38_43 in38 sn43 3183.098862
Rwneg38_44 in38 sn44 3183.098862
Rwneg38_45 in38 sn45 3183.098862
Rwneg38_46 in38 sn46 11140.846016
Rwneg38_47 in38 sn47 11140.846016
Rwneg38_48 in38 sn48 11140.846016
Rwneg38_49 in38 sn49 3183.098862
Rwneg38_50 in38 sn50 11140.846016
Rwneg38_51 in38 sn51 11140.846016
Rwneg38_52 in38 sn52 3183.098862
Rwneg38_53 in38 sn53 11140.846016
Rwneg38_54 in38 sn54 11140.846016
Rwneg38_55 in38 sn55 11140.846016
Rwneg38_56 in38 sn56 11140.846016
Rwneg38_57 in38 sn57 3183.098862
Rwneg38_58 in38 sn58 11140.846016
Rwneg38_59 in38 sn59 3183.098862
Rwneg38_60 in38 sn60 11140.846016
Rwneg38_61 in38 sn61 3183.098862
Rwneg38_62 in38 sn62 11140.846016
Rwneg38_63 in38 sn63 3183.098862
Rwneg38_64 in38 sn64 11140.846016
Rwneg38_65 in38 sn65 3183.098862
Rwneg38_66 in38 sn66 11140.846016
Rwneg38_67 in38 sn67 11140.846016
Rwneg38_68 in38 sn68 11140.846016
Rwneg38_69 in38 sn69 3183.098862
Rwneg38_70 in38 sn70 11140.846016
Rwneg38_71 in38 sn71 11140.846016
Rwneg38_72 in38 sn72 11140.846016
Rwneg38_73 in38 sn73 3183.098862
Rwneg38_74 in38 sn74 11140.846016
Rwneg38_75 in38 sn75 3183.098862
Rwneg38_76 in38 sn76 11140.846016
Rwneg38_77 in38 sn77 3183.098862
Rwneg38_78 in38 sn78 11140.846016
Rwneg38_79 in38 sn79 3183.098862
Rwneg38_80 in38 sn80 3183.098862
Rwneg38_81 in38 sn81 11140.846016
Rwneg38_82 in38 sn82 3183.098862
Rwneg38_83 in38 sn83 3183.098862
Rwneg38_84 in38 sn84 11140.846016
Rwneg38_85 in38 sn85 11140.846016
Rwneg38_86 in38 sn86 11140.846016
Rwneg38_87 in38 sn87 11140.846016
Rwneg38_88 in38 sn88 11140.846016
Rwneg38_89 in38 sn89 3183.098862
Rwneg38_90 in38 sn90 3183.098862
Rwneg38_91 in38 sn91 3183.098862
Rwneg38_92 in38 sn92 11140.846016
Rwneg38_93 in38 sn93 11140.846016
Rwneg38_94 in38 sn94 11140.846016
Rwneg38_95 in38 sn95 3183.098862
Rwneg38_96 in38 sn96 3183.098862
Rwneg38_97 in38 sn97 3183.098862
Rwneg38_98 in38 sn98 11140.846016
Rwneg38_99 in38 sn99 11140.846016
Rwneg38_100 in38 sn100 11140.846016
Rwneg39_1 in39 sn1 3183.098862
Rwneg39_2 in39 sn2 11140.846016
Rwneg39_3 in39 sn3 3183.098862
Rwneg39_4 in39 sn4 11140.846016
Rwneg39_5 in39 sn5 11140.846016
Rwneg39_6 in39 sn6 11140.846016
Rwneg39_7 in39 sn7 11140.846016
Rwneg39_8 in39 sn8 3183.098862
Rwneg39_9 in39 sn9 11140.846016
Rwneg39_10 in39 sn10 11140.846016
Rwneg39_11 in39 sn11 3183.098862
Rwneg39_12 in39 sn12 11140.846016
Rwneg39_13 in39 sn13 11140.846016
Rwneg39_14 in39 sn14 11140.846016
Rwneg39_15 in39 sn15 3183.098862
Rwneg39_16 in39 sn16 11140.846016
Rwneg39_17 in39 sn17 11140.846016
Rwneg39_18 in39 sn18 11140.846016
Rwneg39_19 in39 sn19 11140.846016
Rwneg39_20 in39 sn20 3183.098862
Rwneg39_21 in39 sn21 11140.846016
Rwneg39_22 in39 sn22 11140.846016
Rwneg39_23 in39 sn23 3183.098862
Rwneg39_24 in39 sn24 11140.846016
Rwneg39_25 in39 sn25 3183.098862
Rwneg39_26 in39 sn26 11140.846016
Rwneg39_27 in39 sn27 3183.098862
Rwneg39_28 in39 sn28 3183.098862
Rwneg39_29 in39 sn29 3183.098862
Rwneg39_30 in39 sn30 11140.846016
Rwneg39_31 in39 sn31 11140.846016
Rwneg39_32 in39 sn32 11140.846016
Rwneg39_33 in39 sn33 11140.846016
Rwneg39_34 in39 sn34 11140.846016
Rwneg39_35 in39 sn35 3183.098862
Rwneg39_36 in39 sn36 3183.098862
Rwneg39_37 in39 sn37 11140.846016
Rwneg39_38 in39 sn38 3183.098862
Rwneg39_39 in39 sn39 11140.846016
Rwneg39_40 in39 sn40 11140.846016
Rwneg39_41 in39 sn41 11140.846016
Rwneg39_42 in39 sn42 11140.846016
Rwneg39_43 in39 sn43 3183.098862
Rwneg39_44 in39 sn44 3183.098862
Rwneg39_45 in39 sn45 3183.098862
Rwneg39_46 in39 sn46 11140.846016
Rwneg39_47 in39 sn47 11140.846016
Rwneg39_48 in39 sn48 3183.098862
Rwneg39_49 in39 sn49 3183.098862
Rwneg39_50 in39 sn50 11140.846016
Rwneg39_51 in39 sn51 3183.098862
Rwneg39_52 in39 sn52 3183.098862
Rwneg39_53 in39 sn53 11140.846016
Rwneg39_54 in39 sn54 11140.846016
Rwneg39_55 in39 sn55 3183.098862
Rwneg39_56 in39 sn56 11140.846016
Rwneg39_57 in39 sn57 3183.098862
Rwneg39_58 in39 sn58 11140.846016
Rwneg39_59 in39 sn59 3183.098862
Rwneg39_60 in39 sn60 3183.098862
Rwneg39_61 in39 sn61 11140.846016
Rwneg39_62 in39 sn62 11140.846016
Rwneg39_63 in39 sn63 11140.846016
Rwneg39_64 in39 sn64 11140.846016
Rwneg39_65 in39 sn65 3183.098862
Rwneg39_66 in39 sn66 11140.846016
Rwneg39_67 in39 sn67 11140.846016
Rwneg39_68 in39 sn68 3183.098862
Rwneg39_69 in39 sn69 11140.846016
Rwneg39_70 in39 sn70 11140.846016
Rwneg39_71 in39 sn71 3183.098862
Rwneg39_72 in39 sn72 11140.846016
Rwneg39_73 in39 sn73 3183.098862
Rwneg39_74 in39 sn74 11140.846016
Rwneg39_75 in39 sn75 11140.846016
Rwneg39_76 in39 sn76 11140.846016
Rwneg39_77 in39 sn77 3183.098862
Rwneg39_78 in39 sn78 11140.846016
Rwneg39_79 in39 sn79 11140.846016
Rwneg39_80 in39 sn80 11140.846016
Rwneg39_81 in39 sn81 3183.098862
Rwneg39_82 in39 sn82 11140.846016
Rwneg39_83 in39 sn83 3183.098862
Rwneg39_84 in39 sn84 11140.846016
Rwneg39_85 in39 sn85 3183.098862
Rwneg39_86 in39 sn86 3183.098862
Rwneg39_87 in39 sn87 3183.098862
Rwneg39_88 in39 sn88 11140.846016
Rwneg39_89 in39 sn89 3183.098862
Rwneg39_90 in39 sn90 11140.846016
Rwneg39_91 in39 sn91 11140.846016
Rwneg39_92 in39 sn92 3183.098862
Rwneg39_93 in39 sn93 11140.846016
Rwneg39_94 in39 sn94 11140.846016
Rwneg39_95 in39 sn95 3183.098862
Rwneg39_96 in39 sn96 11140.846016
Rwneg39_97 in39 sn97 11140.846016
Rwneg39_98 in39 sn98 11140.846016
Rwneg39_99 in39 sn99 11140.846016
Rwneg39_100 in39 sn100 11140.846016
Rwneg40_1 in40 sn1 3183.098862
Rwneg40_2 in40 sn2 11140.846016
Rwneg40_3 in40 sn3 11140.846016
Rwneg40_4 in40 sn4 11140.846016
Rwneg40_5 in40 sn5 3183.098862
Rwneg40_6 in40 sn6 3183.098862
Rwneg40_7 in40 sn7 11140.846016
Rwneg40_8 in40 sn8 11140.846016
Rwneg40_9 in40 sn9 3183.098862
Rwneg40_10 in40 sn10 11140.846016
Rwneg40_11 in40 sn11 11140.846016
Rwneg40_12 in40 sn12 3183.098862
Rwneg40_13 in40 sn13 11140.846016
Rwneg40_14 in40 sn14 11140.846016
Rwneg40_15 in40 sn15 3183.098862
Rwneg40_16 in40 sn16 11140.846016
Rwneg40_17 in40 sn17 3183.098862
Rwneg40_18 in40 sn18 3183.098862
Rwneg40_19 in40 sn19 11140.846016
Rwneg40_20 in40 sn20 11140.846016
Rwneg40_21 in40 sn21 3183.098862
Rwneg40_22 in40 sn22 11140.846016
Rwneg40_23 in40 sn23 11140.846016
Rwneg40_24 in40 sn24 3183.098862
Rwneg40_25 in40 sn25 11140.846016
Rwneg40_26 in40 sn26 11140.846016
Rwneg40_27 in40 sn27 11140.846016
Rwneg40_28 in40 sn28 11140.846016
Rwneg40_29 in40 sn29 3183.098862
Rwneg40_30 in40 sn30 11140.846016
Rwneg40_31 in40 sn31 3183.098862
Rwneg40_32 in40 sn32 3183.098862
Rwneg40_33 in40 sn33 3183.098862
Rwneg40_34 in40 sn34 11140.846016
Rwneg40_35 in40 sn35 3183.098862
Rwneg40_36 in40 sn36 11140.846016
Rwneg40_37 in40 sn37 3183.098862
Rwneg40_38 in40 sn38 3183.098862
Rwneg40_39 in40 sn39 11140.846016
Rwneg40_40 in40 sn40 11140.846016
Rwneg40_41 in40 sn41 11140.846016
Rwneg40_42 in40 sn42 11140.846016
Rwneg40_43 in40 sn43 3183.098862
Rwneg40_44 in40 sn44 11140.846016
Rwneg40_45 in40 sn45 3183.098862
Rwneg40_46 in40 sn46 11140.846016
Rwneg40_47 in40 sn47 11140.846016
Rwneg40_48 in40 sn48 11140.846016
Rwneg40_49 in40 sn49 3183.098862
Rwneg40_50 in40 sn50 11140.846016
Rwneg40_51 in40 sn51 11140.846016
Rwneg40_52 in40 sn52 11140.846016
Rwneg40_53 in40 sn53 3183.098862
Rwneg40_54 in40 sn54 3183.098862
Rwneg40_55 in40 sn55 11140.846016
Rwneg40_56 in40 sn56 11140.846016
Rwneg40_57 in40 sn57 11140.846016
Rwneg40_58 in40 sn58 11140.846016
Rwneg40_59 in40 sn59 3183.098862
Rwneg40_60 in40 sn60 11140.846016
Rwneg40_61 in40 sn61 3183.098862
Rwneg40_62 in40 sn62 11140.846016
Rwneg40_63 in40 sn63 11140.846016
Rwneg40_64 in40 sn64 11140.846016
Rwneg40_65 in40 sn65 3183.098862
Rwneg40_66 in40 sn66 3183.098862
Rwneg40_67 in40 sn67 11140.846016
Rwneg40_68 in40 sn68 11140.846016
Rwneg40_69 in40 sn69 11140.846016
Rwneg40_70 in40 sn70 11140.846016
Rwneg40_71 in40 sn71 3183.098862
Rwneg40_72 in40 sn72 11140.846016
Rwneg40_73 in40 sn73 3183.098862
Rwneg40_74 in40 sn74 3183.098862
Rwneg40_75 in40 sn75 3183.098862
Rwneg40_76 in40 sn76 11140.846016
Rwneg40_77 in40 sn77 3183.098862
Rwneg40_78 in40 sn78 11140.846016
Rwneg40_79 in40 sn79 11140.846016
Rwneg40_80 in40 sn80 11140.846016
Rwneg40_81 in40 sn81 3183.098862
Rwneg40_82 in40 sn82 11140.846016
Rwneg40_83 in40 sn83 11140.846016
Rwneg40_84 in40 sn84 11140.846016
Rwneg40_85 in40 sn85 11140.846016
Rwneg40_86 in40 sn86 11140.846016
Rwneg40_87 in40 sn87 11140.846016
Rwneg40_88 in40 sn88 3183.098862
Rwneg40_89 in40 sn89 11140.846016
Rwneg40_90 in40 sn90 11140.846016
Rwneg40_91 in40 sn91 3183.098862
Rwneg40_92 in40 sn92 3183.098862
Rwneg40_93 in40 sn93 3183.098862
Rwneg40_94 in40 sn94 11140.846016
Rwneg40_95 in40 sn95 11140.846016
Rwneg40_96 in40 sn96 11140.846016
Rwneg40_97 in40 sn97 3183.098862
Rwneg40_98 in40 sn98 11140.846016
Rwneg40_99 in40 sn99 11140.846016
Rwneg40_100 in40 sn100 11140.846016
Rwneg41_1 in41 sn1 3183.098862
Rwneg41_2 in41 sn2 11140.846016
Rwneg41_3 in41 sn3 11140.846016
Rwneg41_4 in41 sn4 3183.098862
Rwneg41_5 in41 sn5 11140.846016
Rwneg41_6 in41 sn6 11140.846016
Rwneg41_7 in41 sn7 3183.098862
Rwneg41_8 in41 sn8 11140.846016
Rwneg41_9 in41 sn9 3183.098862
Rwneg41_10 in41 sn10 3183.098862
Rwneg41_11 in41 sn11 11140.846016
Rwneg41_12 in41 sn12 11140.846016
Rwneg41_13 in41 sn13 3183.098862
Rwneg41_14 in41 sn14 11140.846016
Rwneg41_15 in41 sn15 11140.846016
Rwneg41_16 in41 sn16 3183.098862
Rwneg41_17 in41 sn17 3183.098862
Rwneg41_18 in41 sn18 3183.098862
Rwneg41_19 in41 sn19 11140.846016
Rwneg41_20 in41 sn20 3183.098862
Rwneg41_21 in41 sn21 11140.846016
Rwneg41_22 in41 sn22 11140.846016
Rwneg41_23 in41 sn23 11140.846016
Rwneg41_24 in41 sn24 3183.098862
Rwneg41_25 in41 sn25 11140.846016
Rwneg41_26 in41 sn26 3183.098862
Rwneg41_27 in41 sn27 3183.098862
Rwneg41_28 in41 sn28 11140.846016
Rwneg41_29 in41 sn29 11140.846016
Rwneg41_30 in41 sn30 3183.098862
Rwneg41_31 in41 sn31 11140.846016
Rwneg41_32 in41 sn32 3183.098862
Rwneg41_33 in41 sn33 11140.846016
Rwneg41_34 in41 sn34 11140.846016
Rwneg41_35 in41 sn35 3183.098862
Rwneg41_36 in41 sn36 11140.846016
Rwneg41_37 in41 sn37 11140.846016
Rwneg41_38 in41 sn38 11140.846016
Rwneg41_39 in41 sn39 11140.846016
Rwneg41_40 in41 sn40 11140.846016
Rwneg41_41 in41 sn41 11140.846016
Rwneg41_42 in41 sn42 11140.846016
Rwneg41_43 in41 sn43 3183.098862
Rwneg41_44 in41 sn44 11140.846016
Rwneg41_45 in41 sn45 11140.846016
Rwneg41_46 in41 sn46 3183.098862
Rwneg41_47 in41 sn47 11140.846016
Rwneg41_48 in41 sn48 11140.846016
Rwneg41_49 in41 sn49 3183.098862
Rwneg41_50 in41 sn50 3183.098862
Rwneg41_51 in41 sn51 3183.098862
Rwneg41_52 in41 sn52 3183.098862
Rwneg41_53 in41 sn53 3183.098862
Rwneg41_54 in41 sn54 11140.846016
Rwneg41_55 in41 sn55 11140.846016
Rwneg41_56 in41 sn56 3183.098862
Rwneg41_57 in41 sn57 3183.098862
Rwneg41_58 in41 sn58 3183.098862
Rwneg41_59 in41 sn59 3183.098862
Rwneg41_60 in41 sn60 11140.846016
Rwneg41_61 in41 sn61 3183.098862
Rwneg41_62 in41 sn62 3183.098862
Rwneg41_63 in41 sn63 11140.846016
Rwneg41_64 in41 sn64 11140.846016
Rwneg41_65 in41 sn65 3183.098862
Rwneg41_66 in41 sn66 11140.846016
Rwneg41_67 in41 sn67 11140.846016
Rwneg41_68 in41 sn68 3183.098862
Rwneg41_69 in41 sn69 3183.098862
Rwneg41_70 in41 sn70 11140.846016
Rwneg41_71 in41 sn71 11140.846016
Rwneg41_72 in41 sn72 11140.846016
Rwneg41_73 in41 sn73 3183.098862
Rwneg41_74 in41 sn74 3183.098862
Rwneg41_75 in41 sn75 3183.098862
Rwneg41_76 in41 sn76 11140.846016
Rwneg41_77 in41 sn77 3183.098862
Rwneg41_78 in41 sn78 3183.098862
Rwneg41_79 in41 sn79 3183.098862
Rwneg41_80 in41 sn80 3183.098862
Rwneg41_81 in41 sn81 3183.098862
Rwneg41_82 in41 sn82 11140.846016
Rwneg41_83 in41 sn83 3183.098862
Rwneg41_84 in41 sn84 3183.098862
Rwneg41_85 in41 sn85 11140.846016
Rwneg41_86 in41 sn86 11140.846016
Rwneg41_87 in41 sn87 11140.846016
Rwneg41_88 in41 sn88 3183.098862
Rwneg41_89 in41 sn89 11140.846016
Rwneg41_90 in41 sn90 11140.846016
Rwneg41_91 in41 sn91 3183.098862
Rwneg41_92 in41 sn92 11140.846016
Rwneg41_93 in41 sn93 11140.846016
Rwneg41_94 in41 sn94 11140.846016
Rwneg41_95 in41 sn95 3183.098862
Rwneg41_96 in41 sn96 11140.846016
Rwneg41_97 in41 sn97 3183.098862
Rwneg41_98 in41 sn98 11140.846016
Rwneg41_99 in41 sn99 11140.846016
Rwneg41_100 in41 sn100 3183.098862
Rwneg42_1 in42 sn1 11140.846016
Rwneg42_2 in42 sn2 11140.846016
Rwneg42_3 in42 sn3 3183.098862
Rwneg42_4 in42 sn4 11140.846016
Rwneg42_5 in42 sn5 11140.846016
Rwneg42_6 in42 sn6 3183.098862
Rwneg42_7 in42 sn7 3183.098862
Rwneg42_8 in42 sn8 11140.846016
Rwneg42_9 in42 sn9 11140.846016
Rwneg42_10 in42 sn10 11140.846016
Rwneg42_11 in42 sn11 3183.098862
Rwneg42_12 in42 sn12 3183.098862
Rwneg42_13 in42 sn13 3183.098862
Rwneg42_14 in42 sn14 3183.098862
Rwneg42_15 in42 sn15 11140.846016
Rwneg42_16 in42 sn16 3183.098862
Rwneg42_17 in42 sn17 3183.098862
Rwneg42_18 in42 sn18 11140.846016
Rwneg42_19 in42 sn19 11140.846016
Rwneg42_20 in42 sn20 11140.846016
Rwneg42_21 in42 sn21 3183.098862
Rwneg42_22 in42 sn22 3183.098862
Rwneg42_23 in42 sn23 3183.098862
Rwneg42_24 in42 sn24 11140.846016
Rwneg42_25 in42 sn25 3183.098862
Rwneg42_26 in42 sn26 3183.098862
Rwneg42_27 in42 sn27 3183.098862
Rwneg42_28 in42 sn28 3183.098862
Rwneg42_29 in42 sn29 3183.098862
Rwneg42_30 in42 sn30 11140.846016
Rwneg42_31 in42 sn31 11140.846016
Rwneg42_32 in42 sn32 11140.846016
Rwneg42_33 in42 sn33 3183.098862
Rwneg42_34 in42 sn34 3183.098862
Rwneg42_35 in42 sn35 11140.846016
Rwneg42_36 in42 sn36 11140.846016
Rwneg42_37 in42 sn37 11140.846016
Rwneg42_38 in42 sn38 11140.846016
Rwneg42_39 in42 sn39 11140.846016
Rwneg42_40 in42 sn40 11140.846016
Rwneg42_41 in42 sn41 11140.846016
Rwneg42_42 in42 sn42 11140.846016
Rwneg42_43 in42 sn43 3183.098862
Rwneg42_44 in42 sn44 3183.098862
Rwneg42_45 in42 sn45 11140.846016
Rwneg42_46 in42 sn46 3183.098862
Rwneg42_47 in42 sn47 11140.846016
Rwneg42_48 in42 sn48 3183.098862
Rwneg42_49 in42 sn49 3183.098862
Rwneg42_50 in42 sn50 11140.846016
Rwneg42_51 in42 sn51 11140.846016
Rwneg42_52 in42 sn52 11140.846016
Rwneg42_53 in42 sn53 3183.098862
Rwneg42_54 in42 sn54 11140.846016
Rwneg42_55 in42 sn55 11140.846016
Rwneg42_56 in42 sn56 11140.846016
Rwneg42_57 in42 sn57 3183.098862
Rwneg42_58 in42 sn58 3183.098862
Rwneg42_59 in42 sn59 3183.098862
Rwneg42_60 in42 sn60 11140.846016
Rwneg42_61 in42 sn61 11140.846016
Rwneg42_62 in42 sn62 3183.098862
Rwneg42_63 in42 sn63 3183.098862
Rwneg42_64 in42 sn64 3183.098862
Rwneg42_65 in42 sn65 3183.098862
Rwneg42_66 in42 sn66 3183.098862
Rwneg42_67 in42 sn67 11140.846016
Rwneg42_68 in42 sn68 11140.846016
Rwneg42_69 in42 sn69 3183.098862
Rwneg42_70 in42 sn70 11140.846016
Rwneg42_71 in42 sn71 11140.846016
Rwneg42_72 in42 sn72 11140.846016
Rwneg42_73 in42 sn73 3183.098862
Rwneg42_74 in42 sn74 11140.846016
Rwneg42_75 in42 sn75 3183.098862
Rwneg42_76 in42 sn76 11140.846016
Rwneg42_77 in42 sn77 11140.846016
Rwneg42_78 in42 sn78 11140.846016
Rwneg42_79 in42 sn79 11140.846016
Rwneg42_80 in42 sn80 11140.846016
Rwneg42_81 in42 sn81 3183.098862
Rwneg42_82 in42 sn82 11140.846016
Rwneg42_83 in42 sn83 11140.846016
Rwneg42_84 in42 sn84 3183.098862
Rwneg42_85 in42 sn85 3183.098862
Rwneg42_86 in42 sn86 11140.846016
Rwneg42_87 in42 sn87 11140.846016
Rwneg42_88 in42 sn88 11140.846016
Rwneg42_89 in42 sn89 3183.098862
Rwneg42_90 in42 sn90 3183.098862
Rwneg42_91 in42 sn91 3183.098862
Rwneg42_92 in42 sn92 11140.846016
Rwneg42_93 in42 sn93 11140.846016
Rwneg42_94 in42 sn94 3183.098862
Rwneg42_95 in42 sn95 11140.846016
Rwneg42_96 in42 sn96 11140.846016
Rwneg42_97 in42 sn97 3183.098862
Rwneg42_98 in42 sn98 11140.846016
Rwneg42_99 in42 sn99 11140.846016
Rwneg42_100 in42 sn100 11140.846016
Rwneg43_1 in43 sn1 11140.846016
Rwneg43_2 in43 sn2 11140.846016
Rwneg43_3 in43 sn3 11140.846016
Rwneg43_4 in43 sn4 11140.846016
Rwneg43_5 in43 sn5 3183.098862
Rwneg43_6 in43 sn6 3183.098862
Rwneg43_7 in43 sn7 11140.846016
Rwneg43_8 in43 sn8 3183.098862
Rwneg43_9 in43 sn9 11140.846016
Rwneg43_10 in43 sn10 11140.846016
Rwneg43_11 in43 sn11 11140.846016
Rwneg43_12 in43 sn12 3183.098862
Rwneg43_13 in43 sn13 3183.098862
Rwneg43_14 in43 sn14 11140.846016
Rwneg43_15 in43 sn15 11140.846016
Rwneg43_16 in43 sn16 3183.098862
Rwneg43_17 in43 sn17 3183.098862
Rwneg43_18 in43 sn18 11140.846016
Rwneg43_19 in43 sn19 11140.846016
Rwneg43_20 in43 sn20 3183.098862
Rwneg43_21 in43 sn21 3183.098862
Rwneg43_22 in43 sn22 3183.098862
Rwneg43_23 in43 sn23 3183.098862
Rwneg43_24 in43 sn24 3183.098862
Rwneg43_25 in43 sn25 11140.846016
Rwneg43_26 in43 sn26 11140.846016
Rwneg43_27 in43 sn27 11140.846016
Rwneg43_28 in43 sn28 11140.846016
Rwneg43_29 in43 sn29 3183.098862
Rwneg43_30 in43 sn30 11140.846016
Rwneg43_31 in43 sn31 11140.846016
Rwneg43_32 in43 sn32 3183.098862
Rwneg43_33 in43 sn33 3183.098862
Rwneg43_34 in43 sn34 11140.846016
Rwneg43_35 in43 sn35 11140.846016
Rwneg43_36 in43 sn36 11140.846016
Rwneg43_37 in43 sn37 3183.098862
Rwneg43_38 in43 sn38 3183.098862
Rwneg43_39 in43 sn39 3183.098862
Rwneg43_40 in43 sn40 11140.846016
Rwneg43_41 in43 sn41 3183.098862
Rwneg43_42 in43 sn42 11140.846016
Rwneg43_43 in43 sn43 3183.098862
Rwneg43_44 in43 sn44 3183.098862
Rwneg43_45 in43 sn45 3183.098862
Rwneg43_46 in43 sn46 11140.846016
Rwneg43_47 in43 sn47 3183.098862
Rwneg43_48 in43 sn48 11140.846016
Rwneg43_49 in43 sn49 11140.846016
Rwneg43_50 in43 sn50 11140.846016
Rwneg43_51 in43 sn51 11140.846016
Rwneg43_52 in43 sn52 3183.098862
Rwneg43_53 in43 sn53 3183.098862
Rwneg43_54 in43 sn54 3183.098862
Rwneg43_55 in43 sn55 3183.098862
Rwneg43_56 in43 sn56 3183.098862
Rwneg43_57 in43 sn57 3183.098862
Rwneg43_58 in43 sn58 11140.846016
Rwneg43_59 in43 sn59 3183.098862
Rwneg43_60 in43 sn60 3183.098862
Rwneg43_61 in43 sn61 11140.846016
Rwneg43_62 in43 sn62 11140.846016
Rwneg43_63 in43 sn63 3183.098862
Rwneg43_64 in43 sn64 3183.098862
Rwneg43_65 in43 sn65 3183.098862
Rwneg43_66 in43 sn66 11140.846016
Rwneg43_67 in43 sn67 3183.098862
Rwneg43_68 in43 sn68 3183.098862
Rwneg43_69 in43 sn69 11140.846016
Rwneg43_70 in43 sn70 3183.098862
Rwneg43_71 in43 sn71 3183.098862
Rwneg43_72 in43 sn72 11140.846016
Rwneg43_73 in43 sn73 3183.098862
Rwneg43_74 in43 sn74 11140.846016
Rwneg43_75 in43 sn75 3183.098862
Rwneg43_76 in43 sn76 3183.098862
Rwneg43_77 in43 sn77 3183.098862
Rwneg43_78 in43 sn78 11140.846016
Rwneg43_79 in43 sn79 3183.098862
Rwneg43_80 in43 sn80 11140.846016
Rwneg43_81 in43 sn81 11140.846016
Rwneg43_82 in43 sn82 11140.846016
Rwneg43_83 in43 sn83 3183.098862
Rwneg43_84 in43 sn84 3183.098862
Rwneg43_85 in43 sn85 11140.846016
Rwneg43_86 in43 sn86 11140.846016
Rwneg43_87 in43 sn87 3183.098862
Rwneg43_88 in43 sn88 11140.846016
Rwneg43_89 in43 sn89 3183.098862
Rwneg43_90 in43 sn90 11140.846016
Rwneg43_91 in43 sn91 11140.846016
Rwneg43_92 in43 sn92 3183.098862
Rwneg43_93 in43 sn93 3183.098862
Rwneg43_94 in43 sn94 11140.846016
Rwneg43_95 in43 sn95 3183.098862
Rwneg43_96 in43 sn96 3183.098862
Rwneg43_97 in43 sn97 11140.846016
Rwneg43_98 in43 sn98 11140.846016
Rwneg43_99 in43 sn99 3183.098862
Rwneg43_100 in43 sn100 3183.098862
Rwneg44_1 in44 sn1 11140.846016
Rwneg44_2 in44 sn2 11140.846016
Rwneg44_3 in44 sn3 3183.098862
Rwneg44_4 in44 sn4 11140.846016
Rwneg44_5 in44 sn5 3183.098862
Rwneg44_6 in44 sn6 11140.846016
Rwneg44_7 in44 sn7 11140.846016
Rwneg44_8 in44 sn8 3183.098862
Rwneg44_9 in44 sn9 3183.098862
Rwneg44_10 in44 sn10 11140.846016
Rwneg44_11 in44 sn11 3183.098862
Rwneg44_12 in44 sn12 3183.098862
Rwneg44_13 in44 sn13 11140.846016
Rwneg44_14 in44 sn14 11140.846016
Rwneg44_15 in44 sn15 11140.846016
Rwneg44_16 in44 sn16 3183.098862
Rwneg44_17 in44 sn17 11140.846016
Rwneg44_18 in44 sn18 11140.846016
Rwneg44_19 in44 sn19 3183.098862
Rwneg44_20 in44 sn20 11140.846016
Rwneg44_21 in44 sn21 3183.098862
Rwneg44_22 in44 sn22 11140.846016
Rwneg44_23 in44 sn23 11140.846016
Rwneg44_24 in44 sn24 3183.098862
Rwneg44_25 in44 sn25 3183.098862
Rwneg44_26 in44 sn26 11140.846016
Rwneg44_27 in44 sn27 3183.098862
Rwneg44_28 in44 sn28 3183.098862
Rwneg44_29 in44 sn29 3183.098862
Rwneg44_30 in44 sn30 11140.846016
Rwneg44_31 in44 sn31 3183.098862
Rwneg44_32 in44 sn32 3183.098862
Rwneg44_33 in44 sn33 11140.846016
Rwneg44_34 in44 sn34 11140.846016
Rwneg44_35 in44 sn35 3183.098862
Rwneg44_36 in44 sn36 11140.846016
Rwneg44_37 in44 sn37 3183.098862
Rwneg44_38 in44 sn38 3183.098862
Rwneg44_39 in44 sn39 3183.098862
Rwneg44_40 in44 sn40 11140.846016
Rwneg44_41 in44 sn41 3183.098862
Rwneg44_42 in44 sn42 11140.846016
Rwneg44_43 in44 sn43 11140.846016
Rwneg44_44 in44 sn44 3183.098862
Rwneg44_45 in44 sn45 3183.098862
Rwneg44_46 in44 sn46 11140.846016
Rwneg44_47 in44 sn47 3183.098862
Rwneg44_48 in44 sn48 3183.098862
Rwneg44_49 in44 sn49 11140.846016
Rwneg44_50 in44 sn50 3183.098862
Rwneg44_51 in44 sn51 3183.098862
Rwneg44_52 in44 sn52 11140.846016
Rwneg44_53 in44 sn53 3183.098862
Rwneg44_54 in44 sn54 3183.098862
Rwneg44_55 in44 sn55 11140.846016
Rwneg44_56 in44 sn56 3183.098862
Rwneg44_57 in44 sn57 11140.846016
Rwneg44_58 in44 sn58 11140.846016
Rwneg44_59 in44 sn59 3183.098862
Rwneg44_60 in44 sn60 11140.846016
Rwneg44_61 in44 sn61 11140.846016
Rwneg44_62 in44 sn62 11140.846016
Rwneg44_63 in44 sn63 11140.846016
Rwneg44_64 in44 sn64 3183.098862
Rwneg44_65 in44 sn65 11140.846016
Rwneg44_66 in44 sn66 3183.098862
Rwneg44_67 in44 sn67 3183.098862
Rwneg44_68 in44 sn68 11140.846016
Rwneg44_69 in44 sn69 3183.098862
Rwneg44_70 in44 sn70 3183.098862
Rwneg44_71 in44 sn71 11140.846016
Rwneg44_72 in44 sn72 11140.846016
Rwneg44_73 in44 sn73 11140.846016
Rwneg44_74 in44 sn74 11140.846016
Rwneg44_75 in44 sn75 3183.098862
Rwneg44_76 in44 sn76 11140.846016
Rwneg44_77 in44 sn77 3183.098862
Rwneg44_78 in44 sn78 11140.846016
Rwneg44_79 in44 sn79 3183.098862
Rwneg44_80 in44 sn80 3183.098862
Rwneg44_81 in44 sn81 3183.098862
Rwneg44_82 in44 sn82 11140.846016
Rwneg44_83 in44 sn83 11140.846016
Rwneg44_84 in44 sn84 11140.846016
Rwneg44_85 in44 sn85 3183.098862
Rwneg44_86 in44 sn86 3183.098862
Rwneg44_87 in44 sn87 11140.846016
Rwneg44_88 in44 sn88 11140.846016
Rwneg44_89 in44 sn89 3183.098862
Rwneg44_90 in44 sn90 11140.846016
Rwneg44_91 in44 sn91 11140.846016
Rwneg44_92 in44 sn92 3183.098862
Rwneg44_93 in44 sn93 3183.098862
Rwneg44_94 in44 sn94 11140.846016
Rwneg44_95 in44 sn95 11140.846016
Rwneg44_96 in44 sn96 3183.098862
Rwneg44_97 in44 sn97 3183.098862
Rwneg44_98 in44 sn98 3183.098862
Rwneg44_99 in44 sn99 3183.098862
Rwneg44_100 in44 sn100 11140.846016
Rwneg45_1 in45 sn1 11140.846016
Rwneg45_2 in45 sn2 3183.098862
Rwneg45_3 in45 sn3 11140.846016
Rwneg45_4 in45 sn4 11140.846016
Rwneg45_5 in45 sn5 11140.846016
Rwneg45_6 in45 sn6 11140.846016
Rwneg45_7 in45 sn7 3183.098862
Rwneg45_8 in45 sn8 11140.846016
Rwneg45_9 in45 sn9 3183.098862
Rwneg45_10 in45 sn10 11140.846016
Rwneg45_11 in45 sn11 11140.846016
Rwneg45_12 in45 sn12 11140.846016
Rwneg45_13 in45 sn13 3183.098862
Rwneg45_14 in45 sn14 3183.098862
Rwneg45_15 in45 sn15 3183.098862
Rwneg45_16 in45 sn16 11140.846016
Rwneg45_17 in45 sn17 11140.846016
Rwneg45_18 in45 sn18 3183.098862
Rwneg45_19 in45 sn19 11140.846016
Rwneg45_20 in45 sn20 11140.846016
Rwneg45_21 in45 sn21 3183.098862
Rwneg45_22 in45 sn22 11140.846016
Rwneg45_23 in45 sn23 3183.098862
Rwneg45_24 in45 sn24 11140.846016
Rwneg45_25 in45 sn25 3183.098862
Rwneg45_26 in45 sn26 11140.846016
Rwneg45_27 in45 sn27 11140.846016
Rwneg45_28 in45 sn28 11140.846016
Rwneg45_29 in45 sn29 3183.098862
Rwneg45_30 in45 sn30 11140.846016
Rwneg45_31 in45 sn31 11140.846016
Rwneg45_32 in45 sn32 11140.846016
Rwneg45_33 in45 sn33 11140.846016
Rwneg45_34 in45 sn34 11140.846016
Rwneg45_35 in45 sn35 11140.846016
Rwneg45_36 in45 sn36 11140.846016
Rwneg45_37 in45 sn37 11140.846016
Rwneg45_38 in45 sn38 11140.846016
Rwneg45_39 in45 sn39 3183.098862
Rwneg45_40 in45 sn40 3183.098862
Rwneg45_41 in45 sn41 3183.098862
Rwneg45_42 in45 sn42 11140.846016
Rwneg45_43 in45 sn43 3183.098862
Rwneg45_44 in45 sn44 3183.098862
Rwneg45_45 in45 sn45 3183.098862
Rwneg45_46 in45 sn46 11140.846016
Rwneg45_47 in45 sn47 11140.846016
Rwneg45_48 in45 sn48 11140.846016
Rwneg45_49 in45 sn49 3183.098862
Rwneg45_50 in45 sn50 3183.098862
Rwneg45_51 in45 sn51 3183.098862
Rwneg45_52 in45 sn52 3183.098862
Rwneg45_53 in45 sn53 3183.098862
Rwneg45_54 in45 sn54 3183.098862
Rwneg45_55 in45 sn55 3183.098862
Rwneg45_56 in45 sn56 11140.846016
Rwneg45_57 in45 sn57 11140.846016
Rwneg45_58 in45 sn58 11140.846016
Rwneg45_59 in45 sn59 3183.098862
Rwneg45_60 in45 sn60 11140.846016
Rwneg45_61 in45 sn61 11140.846016
Rwneg45_62 in45 sn62 3183.098862
Rwneg45_63 in45 sn63 11140.846016
Rwneg45_64 in45 sn64 11140.846016
Rwneg45_65 in45 sn65 11140.846016
Rwneg45_66 in45 sn66 3183.098862
Rwneg45_67 in45 sn67 11140.846016
Rwneg45_68 in45 sn68 3183.098862
Rwneg45_69 in45 sn69 3183.098862
Rwneg45_70 in45 sn70 11140.846016
Rwneg45_71 in45 sn71 11140.846016
Rwneg45_72 in45 sn72 11140.846016
Rwneg45_73 in45 sn73 11140.846016
Rwneg45_74 in45 sn74 11140.846016
Rwneg45_75 in45 sn75 11140.846016
Rwneg45_76 in45 sn76 3183.098862
Rwneg45_77 in45 sn77 3183.098862
Rwneg45_78 in45 sn78 3183.098862
Rwneg45_79 in45 sn79 11140.846016
Rwneg45_80 in45 sn80 3183.098862
Rwneg45_81 in45 sn81 11140.846016
Rwneg45_82 in45 sn82 11140.846016
Rwneg45_83 in45 sn83 3183.098862
Rwneg45_84 in45 sn84 3183.098862
Rwneg45_85 in45 sn85 11140.846016
Rwneg45_86 in45 sn86 3183.098862
Rwneg45_87 in45 sn87 11140.846016
Rwneg45_88 in45 sn88 11140.846016
Rwneg45_89 in45 sn89 11140.846016
Rwneg45_90 in45 sn90 11140.846016
Rwneg45_91 in45 sn91 3183.098862
Rwneg45_92 in45 sn92 11140.846016
Rwneg45_93 in45 sn93 3183.098862
Rwneg45_94 in45 sn94 3183.098862
Rwneg45_95 in45 sn95 11140.846016
Rwneg45_96 in45 sn96 11140.846016
Rwneg45_97 in45 sn97 3183.098862
Rwneg45_98 in45 sn98 11140.846016
Rwneg45_99 in45 sn99 11140.846016
Rwneg45_100 in45 sn100 11140.846016
Rwneg46_1 in46 sn1 3183.098862
Rwneg46_2 in46 sn2 11140.846016
Rwneg46_3 in46 sn3 3183.098862
Rwneg46_4 in46 sn4 11140.846016
Rwneg46_5 in46 sn5 11140.846016
Rwneg46_6 in46 sn6 3183.098862
Rwneg46_7 in46 sn7 11140.846016
Rwneg46_8 in46 sn8 3183.098862
Rwneg46_9 in46 sn9 3183.098862
Rwneg46_10 in46 sn10 3183.098862
Rwneg46_11 in46 sn11 3183.098862
Rwneg46_12 in46 sn12 3183.098862
Rwneg46_13 in46 sn13 3183.098862
Rwneg46_14 in46 sn14 11140.846016
Rwneg46_15 in46 sn15 11140.846016
Rwneg46_16 in46 sn16 3183.098862
Rwneg46_17 in46 sn17 11140.846016
Rwneg46_18 in46 sn18 3183.098862
Rwneg46_19 in46 sn19 11140.846016
Rwneg46_20 in46 sn20 3183.098862
Rwneg46_21 in46 sn21 3183.098862
Rwneg46_22 in46 sn22 11140.846016
Rwneg46_23 in46 sn23 11140.846016
Rwneg46_24 in46 sn24 3183.098862
Rwneg46_25 in46 sn25 3183.098862
Rwneg46_26 in46 sn26 11140.846016
Rwneg46_27 in46 sn27 3183.098862
Rwneg46_28 in46 sn28 3183.098862
Rwneg46_29 in46 sn29 11140.846016
Rwneg46_30 in46 sn30 11140.846016
Rwneg46_31 in46 sn31 3183.098862
Rwneg46_32 in46 sn32 11140.846016
Rwneg46_33 in46 sn33 11140.846016
Rwneg46_34 in46 sn34 3183.098862
Rwneg46_35 in46 sn35 3183.098862
Rwneg46_36 in46 sn36 3183.098862
Rwneg46_37 in46 sn37 11140.846016
Rwneg46_38 in46 sn38 3183.098862
Rwneg46_39 in46 sn39 11140.846016
Rwneg46_40 in46 sn40 11140.846016
Rwneg46_41 in46 sn41 3183.098862
Rwneg46_42 in46 sn42 3183.098862
Rwneg46_43 in46 sn43 3183.098862
Rwneg46_44 in46 sn44 3183.098862
Rwneg46_45 in46 sn45 3183.098862
Rwneg46_46 in46 sn46 3183.098862
Rwneg46_47 in46 sn47 11140.846016
Rwneg46_48 in46 sn48 3183.098862
Rwneg46_49 in46 sn49 3183.098862
Rwneg46_50 in46 sn50 3183.098862
Rwneg46_51 in46 sn51 3183.098862
Rwneg46_52 in46 sn52 3183.098862
Rwneg46_53 in46 sn53 11140.846016
Rwneg46_54 in46 sn54 11140.846016
Rwneg46_55 in46 sn55 11140.846016
Rwneg46_56 in46 sn56 3183.098862
Rwneg46_57 in46 sn57 3183.098862
Rwneg46_58 in46 sn58 3183.098862
Rwneg46_59 in46 sn59 11140.846016
Rwneg46_60 in46 sn60 11140.846016
Rwneg46_61 in46 sn61 3183.098862
Rwneg46_62 in46 sn62 3183.098862
Rwneg46_63 in46 sn63 11140.846016
Rwneg46_64 in46 sn64 3183.098862
Rwneg46_65 in46 sn65 3183.098862
Rwneg46_66 in46 sn66 3183.098862
Rwneg46_67 in46 sn67 11140.846016
Rwneg46_68 in46 sn68 3183.098862
Rwneg46_69 in46 sn69 11140.846016
Rwneg46_70 in46 sn70 3183.098862
Rwneg46_71 in46 sn71 3183.098862
Rwneg46_72 in46 sn72 3183.098862
Rwneg46_73 in46 sn73 11140.846016
Rwneg46_74 in46 sn74 3183.098862
Rwneg46_75 in46 sn75 3183.098862
Rwneg46_76 in46 sn76 3183.098862
Rwneg46_77 in46 sn77 11140.846016
Rwneg46_78 in46 sn78 3183.098862
Rwneg46_79 in46 sn79 3183.098862
Rwneg46_80 in46 sn80 3183.098862
Rwneg46_81 in46 sn81 11140.846016
Rwneg46_82 in46 sn82 11140.846016
Rwneg46_83 in46 sn83 11140.846016
Rwneg46_84 in46 sn84 3183.098862
Rwneg46_85 in46 sn85 3183.098862
Rwneg46_86 in46 sn86 3183.098862
Rwneg46_87 in46 sn87 11140.846016
Rwneg46_88 in46 sn88 11140.846016
Rwneg46_89 in46 sn89 3183.098862
Rwneg46_90 in46 sn90 11140.846016
Rwneg46_91 in46 sn91 3183.098862
Rwneg46_92 in46 sn92 11140.846016
Rwneg46_93 in46 sn93 3183.098862
Rwneg46_94 in46 sn94 11140.846016
Rwneg46_95 in46 sn95 11140.846016
Rwneg46_96 in46 sn96 11140.846016
Rwneg46_97 in46 sn97 11140.846016
Rwneg46_98 in46 sn98 11140.846016
Rwneg46_99 in46 sn99 11140.846016
Rwneg46_100 in46 sn100 11140.846016
Rwneg47_1 in47 sn1 11140.846016
Rwneg47_2 in47 sn2 3183.098862
Rwneg47_3 in47 sn3 11140.846016
Rwneg47_4 in47 sn4 11140.846016
Rwneg47_5 in47 sn5 3183.098862
Rwneg47_6 in47 sn6 3183.098862
Rwneg47_7 in47 sn7 11140.846016
Rwneg47_8 in47 sn8 3183.098862
Rwneg47_9 in47 sn9 11140.846016
Rwneg47_10 in47 sn10 3183.098862
Rwneg47_11 in47 sn11 11140.846016
Rwneg47_12 in47 sn12 3183.098862
Rwneg47_13 in47 sn13 11140.846016
Rwneg47_14 in47 sn14 11140.846016
Rwneg47_15 in47 sn15 3183.098862
Rwneg47_16 in47 sn16 3183.098862
Rwneg47_17 in47 sn17 3183.098862
Rwneg47_18 in47 sn18 11140.846016
Rwneg47_19 in47 sn19 11140.846016
Rwneg47_20 in47 sn20 11140.846016
Rwneg47_21 in47 sn21 3183.098862
Rwneg47_22 in47 sn22 3183.098862
Rwneg47_23 in47 sn23 11140.846016
Rwneg47_24 in47 sn24 11140.846016
Rwneg47_25 in47 sn25 11140.846016
Rwneg47_26 in47 sn26 11140.846016
Rwneg47_27 in47 sn27 3183.098862
Rwneg47_28 in47 sn28 3183.098862
Rwneg47_29 in47 sn29 3183.098862
Rwneg47_30 in47 sn30 11140.846016
Rwneg47_31 in47 sn31 11140.846016
Rwneg47_32 in47 sn32 11140.846016
Rwneg47_33 in47 sn33 3183.098862
Rwneg47_34 in47 sn34 11140.846016
Rwneg47_35 in47 sn35 11140.846016
Rwneg47_36 in47 sn36 3183.098862
Rwneg47_37 in47 sn37 3183.098862
Rwneg47_38 in47 sn38 3183.098862
Rwneg47_39 in47 sn39 3183.098862
Rwneg47_40 in47 sn40 11140.846016
Rwneg47_41 in47 sn41 11140.846016
Rwneg47_42 in47 sn42 3183.098862
Rwneg47_43 in47 sn43 11140.846016
Rwneg47_44 in47 sn44 3183.098862
Rwneg47_45 in47 sn45 11140.846016
Rwneg47_46 in47 sn46 11140.846016
Rwneg47_47 in47 sn47 11140.846016
Rwneg47_48 in47 sn48 3183.098862
Rwneg47_49 in47 sn49 3183.098862
Rwneg47_50 in47 sn50 11140.846016
Rwneg47_51 in47 sn51 11140.846016
Rwneg47_52 in47 sn52 11140.846016
Rwneg47_53 in47 sn53 3183.098862
Rwneg47_54 in47 sn54 11140.846016
Rwneg47_55 in47 sn55 11140.846016
Rwneg47_56 in47 sn56 11140.846016
Rwneg47_57 in47 sn57 11140.846016
Rwneg47_58 in47 sn58 11140.846016
Rwneg47_59 in47 sn59 3183.098862
Rwneg47_60 in47 sn60 11140.846016
Rwneg47_61 in47 sn61 3183.098862
Rwneg47_62 in47 sn62 11140.846016
Rwneg47_63 in47 sn63 3183.098862
Rwneg47_64 in47 sn64 11140.846016
Rwneg47_65 in47 sn65 3183.098862
Rwneg47_66 in47 sn66 11140.846016
Rwneg47_67 in47 sn67 11140.846016
Rwneg47_68 in47 sn68 11140.846016
Rwneg47_69 in47 sn69 3183.098862
Rwneg47_70 in47 sn70 11140.846016
Rwneg47_71 in47 sn71 3183.098862
Rwneg47_72 in47 sn72 11140.846016
Rwneg47_73 in47 sn73 11140.846016
Rwneg47_74 in47 sn74 11140.846016
Rwneg47_75 in47 sn75 11140.846016
Rwneg47_76 in47 sn76 3183.098862
Rwneg47_77 in47 sn77 3183.098862
Rwneg47_78 in47 sn78 11140.846016
Rwneg47_79 in47 sn79 11140.846016
Rwneg47_80 in47 sn80 3183.098862
Rwneg47_81 in47 sn81 3183.098862
Rwneg47_82 in47 sn82 11140.846016
Rwneg47_83 in47 sn83 11140.846016
Rwneg47_84 in47 sn84 11140.846016
Rwneg47_85 in47 sn85 3183.098862
Rwneg47_86 in47 sn86 11140.846016
Rwneg47_87 in47 sn87 3183.098862
Rwneg47_88 in47 sn88 11140.846016
Rwneg47_89 in47 sn89 3183.098862
Rwneg47_90 in47 sn90 11140.846016
Rwneg47_91 in47 sn91 11140.846016
Rwneg47_92 in47 sn92 3183.098862
Rwneg47_93 in47 sn93 11140.846016
Rwneg47_94 in47 sn94 3183.098862
Rwneg47_95 in47 sn95 11140.846016
Rwneg47_96 in47 sn96 11140.846016
Rwneg47_97 in47 sn97 3183.098862
Rwneg47_98 in47 sn98 11140.846016
Rwneg47_99 in47 sn99 11140.846016
Rwneg47_100 in47 sn100 11140.846016
Rwneg48_1 in48 sn1 3183.098862
Rwneg48_2 in48 sn2 11140.846016
Rwneg48_3 in48 sn3 3183.098862
Rwneg48_4 in48 sn4 11140.846016
Rwneg48_5 in48 sn5 3183.098862
Rwneg48_6 in48 sn6 11140.846016
Rwneg48_7 in48 sn7 3183.098862
Rwneg48_8 in48 sn8 3183.098862
Rwneg48_9 in48 sn9 11140.846016
Rwneg48_10 in48 sn10 11140.846016
Rwneg48_11 in48 sn11 3183.098862
Rwneg48_12 in48 sn12 11140.846016
Rwneg48_13 in48 sn13 3183.098862
Rwneg48_14 in48 sn14 11140.846016
Rwneg48_15 in48 sn15 11140.846016
Rwneg48_16 in48 sn16 11140.846016
Rwneg48_17 in48 sn17 11140.846016
Rwneg48_18 in48 sn18 3183.098862
Rwneg48_19 in48 sn19 3183.098862
Rwneg48_20 in48 sn20 11140.846016
Rwneg48_21 in48 sn21 3183.098862
Rwneg48_22 in48 sn22 11140.846016
Rwneg48_23 in48 sn23 11140.846016
Rwneg48_24 in48 sn24 3183.098862
Rwneg48_25 in48 sn25 11140.846016
Rwneg48_26 in48 sn26 11140.846016
Rwneg48_27 in48 sn27 3183.098862
Rwneg48_28 in48 sn28 3183.098862
Rwneg48_29 in48 sn29 11140.846016
Rwneg48_30 in48 sn30 11140.846016
Rwneg48_31 in48 sn31 3183.098862
Rwneg48_32 in48 sn32 11140.846016
Rwneg48_33 in48 sn33 11140.846016
Rwneg48_34 in48 sn34 11140.846016
Rwneg48_35 in48 sn35 3183.098862
Rwneg48_36 in48 sn36 11140.846016
Rwneg48_37 in48 sn37 3183.098862
Rwneg48_38 in48 sn38 11140.846016
Rwneg48_39 in48 sn39 11140.846016
Rwneg48_40 in48 sn40 3183.098862
Rwneg48_41 in48 sn41 3183.098862
Rwneg48_42 in48 sn42 11140.846016
Rwneg48_43 in48 sn43 3183.098862
Rwneg48_44 in48 sn44 11140.846016
Rwneg48_45 in48 sn45 11140.846016
Rwneg48_46 in48 sn46 11140.846016
Rwneg48_47 in48 sn47 3183.098862
Rwneg48_48 in48 sn48 11140.846016
Rwneg48_49 in48 sn49 11140.846016
Rwneg48_50 in48 sn50 3183.098862
Rwneg48_51 in48 sn51 3183.098862
Rwneg48_52 in48 sn52 11140.846016
Rwneg48_53 in48 sn53 3183.098862
Rwneg48_54 in48 sn54 3183.098862
Rwneg48_55 in48 sn55 11140.846016
Rwneg48_56 in48 sn56 3183.098862
Rwneg48_57 in48 sn57 3183.098862
Rwneg48_58 in48 sn58 11140.846016
Rwneg48_59 in48 sn59 11140.846016
Rwneg48_60 in48 sn60 3183.098862
Rwneg48_61 in48 sn61 11140.846016
Rwneg48_62 in48 sn62 11140.846016
Rwneg48_63 in48 sn63 3183.098862
Rwneg48_64 in48 sn64 3183.098862
Rwneg48_65 in48 sn65 11140.846016
Rwneg48_66 in48 sn66 11140.846016
Rwneg48_67 in48 sn67 3183.098862
Rwneg48_68 in48 sn68 11140.846016
Rwneg48_69 in48 sn69 3183.098862
Rwneg48_70 in48 sn70 3183.098862
Rwneg48_71 in48 sn71 11140.846016
Rwneg48_72 in48 sn72 3183.098862
Rwneg48_73 in48 sn73 11140.846016
Rwneg48_74 in48 sn74 11140.846016
Rwneg48_75 in48 sn75 11140.846016
Rwneg48_76 in48 sn76 11140.846016
Rwneg48_77 in48 sn77 11140.846016
Rwneg48_78 in48 sn78 3183.098862
Rwneg48_79 in48 sn79 3183.098862
Rwneg48_80 in48 sn80 3183.098862
Rwneg48_81 in48 sn81 11140.846016
Rwneg48_82 in48 sn82 3183.098862
Rwneg48_83 in48 sn83 3183.098862
Rwneg48_84 in48 sn84 11140.846016
Rwneg48_85 in48 sn85 3183.098862
Rwneg48_86 in48 sn86 11140.846016
Rwneg48_87 in48 sn87 11140.846016
Rwneg48_88 in48 sn88 3183.098862
Rwneg48_89 in48 sn89 3183.098862
Rwneg48_90 in48 sn90 11140.846016
Rwneg48_91 in48 sn91 11140.846016
Rwneg48_92 in48 sn92 3183.098862
Rwneg48_93 in48 sn93 11140.846016
Rwneg48_94 in48 sn94 11140.846016
Rwneg48_95 in48 sn95 11140.846016
Rwneg48_96 in48 sn96 3183.098862
Rwneg48_97 in48 sn97 11140.846016
Rwneg48_98 in48 sn98 3183.098862
Rwneg48_99 in48 sn99 3183.098862
Rwneg48_100 in48 sn100 11140.846016
Rwneg49_1 in49 sn1 3183.098862
Rwneg49_2 in49 sn2 3183.098862
Rwneg49_3 in49 sn3 3183.098862
Rwneg49_4 in49 sn4 11140.846016
Rwneg49_5 in49 sn5 3183.098862
Rwneg49_6 in49 sn6 11140.846016
Rwneg49_7 in49 sn7 11140.846016
Rwneg49_8 in49 sn8 3183.098862
Rwneg49_9 in49 sn9 11140.846016
Rwneg49_10 in49 sn10 11140.846016
Rwneg49_11 in49 sn11 3183.098862
Rwneg49_12 in49 sn12 3183.098862
Rwneg49_13 in49 sn13 11140.846016
Rwneg49_14 in49 sn14 11140.846016
Rwneg49_15 in49 sn15 3183.098862
Rwneg49_16 in49 sn16 11140.846016
Rwneg49_17 in49 sn17 3183.098862
Rwneg49_18 in49 sn18 3183.098862
Rwneg49_19 in49 sn19 3183.098862
Rwneg49_20 in49 sn20 3183.098862
Rwneg49_21 in49 sn21 11140.846016
Rwneg49_22 in49 sn22 11140.846016
Rwneg49_23 in49 sn23 11140.846016
Rwneg49_24 in49 sn24 11140.846016
Rwneg49_25 in49 sn25 11140.846016
Rwneg49_26 in49 sn26 11140.846016
Rwneg49_27 in49 sn27 11140.846016
Rwneg49_28 in49 sn28 3183.098862
Rwneg49_29 in49 sn29 11140.846016
Rwneg49_30 in49 sn30 3183.098862
Rwneg49_31 in49 sn31 3183.098862
Rwneg49_32 in49 sn32 3183.098862
Rwneg49_33 in49 sn33 3183.098862
Rwneg49_34 in49 sn34 3183.098862
Rwneg49_35 in49 sn35 11140.846016
Rwneg49_36 in49 sn36 3183.098862
Rwneg49_37 in49 sn37 11140.846016
Rwneg49_38 in49 sn38 11140.846016
Rwneg49_39 in49 sn39 11140.846016
Rwneg49_40 in49 sn40 11140.846016
Rwneg49_41 in49 sn41 11140.846016
Rwneg49_42 in49 sn42 11140.846016
Rwneg49_43 in49 sn43 11140.846016
Rwneg49_44 in49 sn44 3183.098862
Rwneg49_45 in49 sn45 3183.098862
Rwneg49_46 in49 sn46 3183.098862
Rwneg49_47 in49 sn47 3183.098862
Rwneg49_48 in49 sn48 11140.846016
Rwneg49_49 in49 sn49 11140.846016
Rwneg49_50 in49 sn50 3183.098862
Rwneg49_51 in49 sn51 11140.846016
Rwneg49_52 in49 sn52 3183.098862
Rwneg49_53 in49 sn53 11140.846016
Rwneg49_54 in49 sn54 11140.846016
Rwneg49_55 in49 sn55 11140.846016
Rwneg49_56 in49 sn56 11140.846016
Rwneg49_57 in49 sn57 3183.098862
Rwneg49_58 in49 sn58 3183.098862
Rwneg49_59 in49 sn59 11140.846016
Rwneg49_60 in49 sn60 3183.098862
Rwneg49_61 in49 sn61 3183.098862
Rwneg49_62 in49 sn62 3183.098862
Rwneg49_63 in49 sn63 3183.098862
Rwneg49_64 in49 sn64 11140.846016
Rwneg49_65 in49 sn65 3183.098862
Rwneg49_66 in49 sn66 3183.098862
Rwneg49_67 in49 sn67 11140.846016
Rwneg49_68 in49 sn68 11140.846016
Rwneg49_69 in49 sn69 11140.846016
Rwneg49_70 in49 sn70 11140.846016
Rwneg49_71 in49 sn71 3183.098862
Rwneg49_72 in49 sn72 11140.846016
Rwneg49_73 in49 sn73 3183.098862
Rwneg49_74 in49 sn74 11140.846016
Rwneg49_75 in49 sn75 3183.098862
Rwneg49_76 in49 sn76 3183.098862
Rwneg49_77 in49 sn77 3183.098862
Rwneg49_78 in49 sn78 11140.846016
Rwneg49_79 in49 sn79 3183.098862
Rwneg49_80 in49 sn80 11140.846016
Rwneg49_81 in49 sn81 3183.098862
Rwneg49_82 in49 sn82 3183.098862
Rwneg49_83 in49 sn83 3183.098862
Rwneg49_84 in49 sn84 11140.846016
Rwneg49_85 in49 sn85 3183.098862
Rwneg49_86 in49 sn86 3183.098862
Rwneg49_87 in49 sn87 11140.846016
Rwneg49_88 in49 sn88 11140.846016
Rwneg49_89 in49 sn89 3183.098862
Rwneg49_90 in49 sn90 11140.846016
Rwneg49_91 in49 sn91 11140.846016
Rwneg49_92 in49 sn92 11140.846016
Rwneg49_93 in49 sn93 3183.098862
Rwneg49_94 in49 sn94 11140.846016
Rwneg49_95 in49 sn95 11140.846016
Rwneg49_96 in49 sn96 11140.846016
Rwneg49_97 in49 sn97 11140.846016
Rwneg49_98 in49 sn98 3183.098862
Rwneg49_99 in49 sn99 11140.846016
Rwneg49_100 in49 sn100 3183.098862
Rwneg50_1 in50 sn1 11140.846016
Rwneg50_2 in50 sn2 3183.098862
Rwneg50_3 in50 sn3 11140.846016
Rwneg50_4 in50 sn4 11140.846016
Rwneg50_5 in50 sn5 3183.098862
Rwneg50_6 in50 sn6 11140.846016
Rwneg50_7 in50 sn7 3183.098862
Rwneg50_8 in50 sn8 3183.098862
Rwneg50_9 in50 sn9 3183.098862
Rwneg50_10 in50 sn10 11140.846016
Rwneg50_11 in50 sn11 3183.098862
Rwneg50_12 in50 sn12 11140.846016
Rwneg50_13 in50 sn13 3183.098862
Rwneg50_14 in50 sn14 3183.098862
Rwneg50_15 in50 sn15 3183.098862
Rwneg50_16 in50 sn16 11140.846016
Rwneg50_17 in50 sn17 11140.846016
Rwneg50_18 in50 sn18 11140.846016
Rwneg50_19 in50 sn19 11140.846016
Rwneg50_20 in50 sn20 3183.098862
Rwneg50_21 in50 sn21 3183.098862
Rwneg50_22 in50 sn22 3183.098862
Rwneg50_23 in50 sn23 11140.846016
Rwneg50_24 in50 sn24 3183.098862
Rwneg50_25 in50 sn25 11140.846016
Rwneg50_26 in50 sn26 11140.846016
Rwneg50_27 in50 sn27 3183.098862
Rwneg50_28 in50 sn28 11140.846016
Rwneg50_29 in50 sn29 11140.846016
Rwneg50_30 in50 sn30 3183.098862
Rwneg50_31 in50 sn31 3183.098862
Rwneg50_32 in50 sn32 3183.098862
Rwneg50_33 in50 sn33 11140.846016
Rwneg50_34 in50 sn34 3183.098862
Rwneg50_35 in50 sn35 3183.098862
Rwneg50_36 in50 sn36 11140.846016
Rwneg50_37 in50 sn37 3183.098862
Rwneg50_38 in50 sn38 3183.098862
Rwneg50_39 in50 sn39 11140.846016
Rwneg50_40 in50 sn40 11140.846016
Rwneg50_41 in50 sn41 11140.846016
Rwneg50_42 in50 sn42 11140.846016
Rwneg50_43 in50 sn43 3183.098862
Rwneg50_44 in50 sn44 3183.098862
Rwneg50_45 in50 sn45 11140.846016
Rwneg50_46 in50 sn46 3183.098862
Rwneg50_47 in50 sn47 11140.846016
Rwneg50_48 in50 sn48 3183.098862
Rwneg50_49 in50 sn49 3183.098862
Rwneg50_50 in50 sn50 11140.846016
Rwneg50_51 in50 sn51 3183.098862
Rwneg50_52 in50 sn52 11140.846016
Rwneg50_53 in50 sn53 11140.846016
Rwneg50_54 in50 sn54 11140.846016
Rwneg50_55 in50 sn55 3183.098862
Rwneg50_56 in50 sn56 11140.846016
Rwneg50_57 in50 sn57 11140.846016
Rwneg50_58 in50 sn58 11140.846016
Rwneg50_59 in50 sn59 11140.846016
Rwneg50_60 in50 sn60 3183.098862
Rwneg50_61 in50 sn61 11140.846016
Rwneg50_62 in50 sn62 3183.098862
Rwneg50_63 in50 sn63 3183.098862
Rwneg50_64 in50 sn64 11140.846016
Rwneg50_65 in50 sn65 11140.846016
Rwneg50_66 in50 sn66 3183.098862
Rwneg50_67 in50 sn67 11140.846016
Rwneg50_68 in50 sn68 3183.098862
Rwneg50_69 in50 sn69 11140.846016
Rwneg50_70 in50 sn70 11140.846016
Rwneg50_71 in50 sn71 11140.846016
Rwneg50_72 in50 sn72 11140.846016
Rwneg50_73 in50 sn73 3183.098862
Rwneg50_74 in50 sn74 11140.846016
Rwneg50_75 in50 sn75 3183.098862
Rwneg50_76 in50 sn76 11140.846016
Rwneg50_77 in50 sn77 3183.098862
Rwneg50_78 in50 sn78 3183.098862
Rwneg50_79 in50 sn79 11140.846016
Rwneg50_80 in50 sn80 3183.098862
Rwneg50_81 in50 sn81 11140.846016
Rwneg50_82 in50 sn82 3183.098862
Rwneg50_83 in50 sn83 11140.846016
Rwneg50_84 in50 sn84 3183.098862
Rwneg50_85 in50 sn85 3183.098862
Rwneg50_86 in50 sn86 11140.846016
Rwneg50_87 in50 sn87 3183.098862
Rwneg50_88 in50 sn88 3183.098862
Rwneg50_89 in50 sn89 11140.846016
Rwneg50_90 in50 sn90 3183.098862
Rwneg50_91 in50 sn91 3183.098862
Rwneg50_92 in50 sn92 3183.098862
Rwneg50_93 in50 sn93 3183.098862
Rwneg50_94 in50 sn94 3183.098862
Rwneg50_95 in50 sn95 3183.098862
Rwneg50_96 in50 sn96 3183.098862
Rwneg50_97 in50 sn97 11140.846016
Rwneg50_98 in50 sn98 11140.846016
Rwneg50_99 in50 sn99 3183.098862
Rwneg50_100 in50 sn100 11140.846016
Rwneg51_1 in51 sn1 3183.098862
Rwneg51_2 in51 sn2 3183.098862
Rwneg51_3 in51 sn3 3183.098862
Rwneg51_4 in51 sn4 11140.846016
Rwneg51_5 in51 sn5 11140.846016
Rwneg51_6 in51 sn6 3183.098862
Rwneg51_7 in51 sn7 11140.846016
Rwneg51_8 in51 sn8 11140.846016
Rwneg51_9 in51 sn9 11140.846016
Rwneg51_10 in51 sn10 3183.098862
Rwneg51_11 in51 sn11 3183.098862
Rwneg51_12 in51 sn12 11140.846016
Rwneg51_13 in51 sn13 3183.098862
Rwneg51_14 in51 sn14 11140.846016
Rwneg51_15 in51 sn15 11140.846016
Rwneg51_16 in51 sn16 11140.846016
Rwneg51_17 in51 sn17 11140.846016
Rwneg51_18 in51 sn18 11140.846016
Rwneg51_19 in51 sn19 11140.846016
Rwneg51_20 in51 sn20 11140.846016
Rwneg51_21 in51 sn21 3183.098862
Rwneg51_22 in51 sn22 3183.098862
Rwneg51_23 in51 sn23 3183.098862
Rwneg51_24 in51 sn24 11140.846016
Rwneg51_25 in51 sn25 11140.846016
Rwneg51_26 in51 sn26 3183.098862
Rwneg51_27 in51 sn27 3183.098862
Rwneg51_28 in51 sn28 3183.098862
Rwneg51_29 in51 sn29 3183.098862
Rwneg51_30 in51 sn30 11140.846016
Rwneg51_31 in51 sn31 3183.098862
Rwneg51_32 in51 sn32 3183.098862
Rwneg51_33 in51 sn33 3183.098862
Rwneg51_34 in51 sn34 11140.846016
Rwneg51_35 in51 sn35 11140.846016
Rwneg51_36 in51 sn36 11140.846016
Rwneg51_37 in51 sn37 11140.846016
Rwneg51_38 in51 sn38 3183.098862
Rwneg51_39 in51 sn39 3183.098862
Rwneg51_40 in51 sn40 11140.846016
Rwneg51_41 in51 sn41 11140.846016
Rwneg51_42 in51 sn42 11140.846016
Rwneg51_43 in51 sn43 3183.098862
Rwneg51_44 in51 sn44 3183.098862
Rwneg51_45 in51 sn45 3183.098862
Rwneg51_46 in51 sn46 11140.846016
Rwneg51_47 in51 sn47 11140.846016
Rwneg51_48 in51 sn48 3183.098862
Rwneg51_49 in51 sn49 3183.098862
Rwneg51_50 in51 sn50 3183.098862
Rwneg51_51 in51 sn51 11140.846016
Rwneg51_52 in51 sn52 11140.846016
Rwneg51_53 in51 sn53 3183.098862
Rwneg51_54 in51 sn54 3183.098862
Rwneg51_55 in51 sn55 3183.098862
Rwneg51_56 in51 sn56 11140.846016
Rwneg51_57 in51 sn57 11140.846016
Rwneg51_58 in51 sn58 11140.846016
Rwneg51_59 in51 sn59 3183.098862
Rwneg51_60 in51 sn60 11140.846016
Rwneg51_61 in51 sn61 11140.846016
Rwneg51_62 in51 sn62 11140.846016
Rwneg51_63 in51 sn63 11140.846016
Rwneg51_64 in51 sn64 3183.098862
Rwneg51_65 in51 sn65 3183.098862
Rwneg51_66 in51 sn66 3183.098862
Rwneg51_67 in51 sn67 11140.846016
Rwneg51_68 in51 sn68 11140.846016
Rwneg51_69 in51 sn69 3183.098862
Rwneg51_70 in51 sn70 3183.098862
Rwneg51_71 in51 sn71 11140.846016
Rwneg51_72 in51 sn72 11140.846016
Rwneg51_73 in51 sn73 11140.846016
Rwneg51_74 in51 sn74 11140.846016
Rwneg51_75 in51 sn75 3183.098862
Rwneg51_76 in51 sn76 3183.098862
Rwneg51_77 in51 sn77 3183.098862
Rwneg51_78 in51 sn78 11140.846016
Rwneg51_79 in51 sn79 3183.098862
Rwneg51_80 in51 sn80 3183.098862
Rwneg51_81 in51 sn81 11140.846016
Rwneg51_82 in51 sn82 3183.098862
Rwneg51_83 in51 sn83 11140.846016
Rwneg51_84 in51 sn84 11140.846016
Rwneg51_85 in51 sn85 3183.098862
Rwneg51_86 in51 sn86 3183.098862
Rwneg51_87 in51 sn87 11140.846016
Rwneg51_88 in51 sn88 11140.846016
Rwneg51_89 in51 sn89 11140.846016
Rwneg51_90 in51 sn90 3183.098862
Rwneg51_91 in51 sn91 3183.098862
Rwneg51_92 in51 sn92 11140.846016
Rwneg51_93 in51 sn93 3183.098862
Rwneg51_94 in51 sn94 11140.846016
Rwneg51_95 in51 sn95 11140.846016
Rwneg51_96 in51 sn96 11140.846016
Rwneg51_97 in51 sn97 3183.098862
Rwneg51_98 in51 sn98 3183.098862
Rwneg51_99 in51 sn99 11140.846016
Rwneg51_100 in51 sn100 11140.846016
Rwneg52_1 in52 sn1 3183.098862
Rwneg52_2 in52 sn2 3183.098862
Rwneg52_3 in52 sn3 3183.098862
Rwneg52_4 in52 sn4 11140.846016
Rwneg52_5 in52 sn5 11140.846016
Rwneg52_6 in52 sn6 3183.098862
Rwneg52_7 in52 sn7 11140.846016
Rwneg52_8 in52 sn8 11140.846016
Rwneg52_9 in52 sn9 3183.098862
Rwneg52_10 in52 sn10 11140.846016
Rwneg52_11 in52 sn11 3183.098862
Rwneg52_12 in52 sn12 3183.098862
Rwneg52_13 in52 sn13 3183.098862
Rwneg52_14 in52 sn14 3183.098862
Rwneg52_15 in52 sn15 11140.846016
Rwneg52_16 in52 sn16 11140.846016
Rwneg52_17 in52 sn17 3183.098862
Rwneg52_18 in52 sn18 11140.846016
Rwneg52_19 in52 sn19 11140.846016
Rwneg52_20 in52 sn20 11140.846016
Rwneg52_21 in52 sn21 11140.846016
Rwneg52_22 in52 sn22 3183.098862
Rwneg52_23 in52 sn23 3183.098862
Rwneg52_24 in52 sn24 11140.846016
Rwneg52_25 in52 sn25 11140.846016
Rwneg52_26 in52 sn26 11140.846016
Rwneg52_27 in52 sn27 11140.846016
Rwneg52_28 in52 sn28 3183.098862
Rwneg52_29 in52 sn29 3183.098862
Rwneg52_30 in52 sn30 3183.098862
Rwneg52_31 in52 sn31 11140.846016
Rwneg52_32 in52 sn32 11140.846016
Rwneg52_33 in52 sn33 3183.098862
Rwneg52_34 in52 sn34 3183.098862
Rwneg52_35 in52 sn35 3183.098862
Rwneg52_36 in52 sn36 11140.846016
Rwneg52_37 in52 sn37 3183.098862
Rwneg52_38 in52 sn38 3183.098862
Rwneg52_39 in52 sn39 11140.846016
Rwneg52_40 in52 sn40 3183.098862
Rwneg52_41 in52 sn41 3183.098862
Rwneg52_42 in52 sn42 3183.098862
Rwneg52_43 in52 sn43 3183.098862
Rwneg52_44 in52 sn44 11140.846016
Rwneg52_45 in52 sn45 3183.098862
Rwneg52_46 in52 sn46 11140.846016
Rwneg52_47 in52 sn47 11140.846016
Rwneg52_48 in52 sn48 11140.846016
Rwneg52_49 in52 sn49 3183.098862
Rwneg52_50 in52 sn50 11140.846016
Rwneg52_51 in52 sn51 11140.846016
Rwneg52_52 in52 sn52 11140.846016
Rwneg52_53 in52 sn53 3183.098862
Rwneg52_54 in52 sn54 11140.846016
Rwneg52_55 in52 sn55 11140.846016
Rwneg52_56 in52 sn56 3183.098862
Rwneg52_57 in52 sn57 3183.098862
Rwneg52_58 in52 sn58 3183.098862
Rwneg52_59 in52 sn59 3183.098862
Rwneg52_60 in52 sn60 11140.846016
Rwneg52_61 in52 sn61 11140.846016
Rwneg52_62 in52 sn62 11140.846016
Rwneg52_63 in52 sn63 11140.846016
Rwneg52_64 in52 sn64 11140.846016
Rwneg52_65 in52 sn65 11140.846016
Rwneg52_66 in52 sn66 3183.098862
Rwneg52_67 in52 sn67 11140.846016
Rwneg52_68 in52 sn68 11140.846016
Rwneg52_69 in52 sn69 3183.098862
Rwneg52_70 in52 sn70 11140.846016
Rwneg52_71 in52 sn71 3183.098862
Rwneg52_72 in52 sn72 3183.098862
Rwneg52_73 in52 sn73 3183.098862
Rwneg52_74 in52 sn74 3183.098862
Rwneg52_75 in52 sn75 3183.098862
Rwneg52_76 in52 sn76 3183.098862
Rwneg52_77 in52 sn77 11140.846016
Rwneg52_78 in52 sn78 11140.846016
Rwneg52_79 in52 sn79 3183.098862
Rwneg52_80 in52 sn80 11140.846016
Rwneg52_81 in52 sn81 11140.846016
Rwneg52_82 in52 sn82 3183.098862
Rwneg52_83 in52 sn83 11140.846016
Rwneg52_84 in52 sn84 11140.846016
Rwneg52_85 in52 sn85 3183.098862
Rwneg52_86 in52 sn86 3183.098862
Rwneg52_87 in52 sn87 11140.846016
Rwneg52_88 in52 sn88 3183.098862
Rwneg52_89 in52 sn89 3183.098862
Rwneg52_90 in52 sn90 3183.098862
Rwneg52_91 in52 sn91 11140.846016
Rwneg52_92 in52 sn92 3183.098862
Rwneg52_93 in52 sn93 11140.846016
Rwneg52_94 in52 sn94 3183.098862
Rwneg52_95 in52 sn95 3183.098862
Rwneg52_96 in52 sn96 11140.846016
Rwneg52_97 in52 sn97 11140.846016
Rwneg52_98 in52 sn98 11140.846016
Rwneg52_99 in52 sn99 3183.098862
Rwneg52_100 in52 sn100 11140.846016
Rwneg53_1 in53 sn1 3183.098862
Rwneg53_2 in53 sn2 3183.098862
Rwneg53_3 in53 sn3 3183.098862
Rwneg53_4 in53 sn4 11140.846016
Rwneg53_5 in53 sn5 11140.846016
Rwneg53_6 in53 sn6 11140.846016
Rwneg53_7 in53 sn7 11140.846016
Rwneg53_8 in53 sn8 3183.098862
Rwneg53_9 in53 sn9 11140.846016
Rwneg53_10 in53 sn10 11140.846016
Rwneg53_11 in53 sn11 3183.098862
Rwneg53_12 in53 sn12 11140.846016
Rwneg53_13 in53 sn13 11140.846016
Rwneg53_14 in53 sn14 11140.846016
Rwneg53_15 in53 sn15 3183.098862
Rwneg53_16 in53 sn16 11140.846016
Rwneg53_17 in53 sn17 3183.098862
Rwneg53_18 in53 sn18 3183.098862
Rwneg53_19 in53 sn19 3183.098862
Rwneg53_20 in53 sn20 3183.098862
Rwneg53_21 in53 sn21 3183.098862
Rwneg53_22 in53 sn22 3183.098862
Rwneg53_23 in53 sn23 11140.846016
Rwneg53_24 in53 sn24 3183.098862
Rwneg53_25 in53 sn25 11140.846016
Rwneg53_26 in53 sn26 3183.098862
Rwneg53_27 in53 sn27 11140.846016
Rwneg53_28 in53 sn28 3183.098862
Rwneg53_29 in53 sn29 11140.846016
Rwneg53_30 in53 sn30 11140.846016
Rwneg53_31 in53 sn31 3183.098862
Rwneg53_32 in53 sn32 3183.098862
Rwneg53_33 in53 sn33 3183.098862
Rwneg53_34 in53 sn34 3183.098862
Rwneg53_35 in53 sn35 3183.098862
Rwneg53_36 in53 sn36 11140.846016
Rwneg53_37 in53 sn37 11140.846016
Rwneg53_38 in53 sn38 11140.846016
Rwneg53_39 in53 sn39 11140.846016
Rwneg53_40 in53 sn40 3183.098862
Rwneg53_41 in53 sn41 11140.846016
Rwneg53_42 in53 sn42 11140.846016
Rwneg53_43 in53 sn43 3183.098862
Rwneg53_44 in53 sn44 3183.098862
Rwneg53_45 in53 sn45 11140.846016
Rwneg53_46 in53 sn46 3183.098862
Rwneg53_47 in53 sn47 3183.098862
Rwneg53_48 in53 sn48 11140.846016
Rwneg53_49 in53 sn49 3183.098862
Rwneg53_50 in53 sn50 11140.846016
Rwneg53_51 in53 sn51 3183.098862
Rwneg53_52 in53 sn52 3183.098862
Rwneg53_53 in53 sn53 3183.098862
Rwneg53_54 in53 sn54 11140.846016
Rwneg53_55 in53 sn55 11140.846016
Rwneg53_56 in53 sn56 3183.098862
Rwneg53_57 in53 sn57 11140.846016
Rwneg53_58 in53 sn58 11140.846016
Rwneg53_59 in53 sn59 3183.098862
Rwneg53_60 in53 sn60 3183.098862
Rwneg53_61 in53 sn61 11140.846016
Rwneg53_62 in53 sn62 3183.098862
Rwneg53_63 in53 sn63 3183.098862
Rwneg53_64 in53 sn64 11140.846016
Rwneg53_65 in53 sn65 11140.846016
Rwneg53_66 in53 sn66 3183.098862
Rwneg53_67 in53 sn67 3183.098862
Rwneg53_68 in53 sn68 11140.846016
Rwneg53_69 in53 sn69 11140.846016
Rwneg53_70 in53 sn70 11140.846016
Rwneg53_71 in53 sn71 11140.846016
Rwneg53_72 in53 sn72 3183.098862
Rwneg53_73 in53 sn73 11140.846016
Rwneg53_74 in53 sn74 11140.846016
Rwneg53_75 in53 sn75 11140.846016
Rwneg53_76 in53 sn76 3183.098862
Rwneg53_77 in53 sn77 11140.846016
Rwneg53_78 in53 sn78 3183.098862
Rwneg53_79 in53 sn79 3183.098862
Rwneg53_80 in53 sn80 11140.846016
Rwneg53_81 in53 sn81 11140.846016
Rwneg53_82 in53 sn82 3183.098862
Rwneg53_83 in53 sn83 3183.098862
Rwneg53_84 in53 sn84 3183.098862
Rwneg53_85 in53 sn85 3183.098862
Rwneg53_86 in53 sn86 11140.846016
Rwneg53_87 in53 sn87 11140.846016
Rwneg53_88 in53 sn88 3183.098862
Rwneg53_89 in53 sn89 11140.846016
Rwneg53_90 in53 sn90 3183.098862
Rwneg53_91 in53 sn91 11140.846016
Rwneg53_92 in53 sn92 11140.846016
Rwneg53_93 in53 sn93 11140.846016
Rwneg53_94 in53 sn94 3183.098862
Rwneg53_95 in53 sn95 3183.098862
Rwneg53_96 in53 sn96 11140.846016
Rwneg53_97 in53 sn97 11140.846016
Rwneg53_98 in53 sn98 3183.098862
Rwneg53_99 in53 sn99 11140.846016
Rwneg53_100 in53 sn100 11140.846016
Rwneg54_1 in54 sn1 11140.846016
Rwneg54_2 in54 sn2 3183.098862
Rwneg54_3 in54 sn3 3183.098862
Rwneg54_4 in54 sn4 11140.846016
Rwneg54_5 in54 sn5 11140.846016
Rwneg54_6 in54 sn6 11140.846016
Rwneg54_7 in54 sn7 11140.846016
Rwneg54_8 in54 sn8 3183.098862
Rwneg54_9 in54 sn9 3183.098862
Rwneg54_10 in54 sn10 3183.098862
Rwneg54_11 in54 sn11 3183.098862
Rwneg54_12 in54 sn12 11140.846016
Rwneg54_13 in54 sn13 3183.098862
Rwneg54_14 in54 sn14 3183.098862
Rwneg54_15 in54 sn15 3183.098862
Rwneg54_16 in54 sn16 3183.098862
Rwneg54_17 in54 sn17 3183.098862
Rwneg54_18 in54 sn18 3183.098862
Rwneg54_19 in54 sn19 3183.098862
Rwneg54_20 in54 sn20 11140.846016
Rwneg54_21 in54 sn21 11140.846016
Rwneg54_22 in54 sn22 11140.846016
Rwneg54_23 in54 sn23 3183.098862
Rwneg54_24 in54 sn24 3183.098862
Rwneg54_25 in54 sn25 11140.846016
Rwneg54_26 in54 sn26 11140.846016
Rwneg54_27 in54 sn27 3183.098862
Rwneg54_28 in54 sn28 3183.098862
Rwneg54_29 in54 sn29 11140.846016
Rwneg54_30 in54 sn30 11140.846016
Rwneg54_31 in54 sn31 11140.846016
Rwneg54_32 in54 sn32 3183.098862
Rwneg54_33 in54 sn33 11140.846016
Rwneg54_34 in54 sn34 11140.846016
Rwneg54_35 in54 sn35 11140.846016
Rwneg54_36 in54 sn36 11140.846016
Rwneg54_37 in54 sn37 3183.098862
Rwneg54_38 in54 sn38 3183.098862
Rwneg54_39 in54 sn39 3183.098862
Rwneg54_40 in54 sn40 11140.846016
Rwneg54_41 in54 sn41 3183.098862
Rwneg54_42 in54 sn42 3183.098862
Rwneg54_43 in54 sn43 11140.846016
Rwneg54_44 in54 sn44 3183.098862
Rwneg54_45 in54 sn45 3183.098862
Rwneg54_46 in54 sn46 11140.846016
Rwneg54_47 in54 sn47 11140.846016
Rwneg54_48 in54 sn48 11140.846016
Rwneg54_49 in54 sn49 11140.846016
Rwneg54_50 in54 sn50 3183.098862
Rwneg54_51 in54 sn51 11140.846016
Rwneg54_52 in54 sn52 11140.846016
Rwneg54_53 in54 sn53 3183.098862
Rwneg54_54 in54 sn54 11140.846016
Rwneg54_55 in54 sn55 3183.098862
Rwneg54_56 in54 sn56 3183.098862
Rwneg54_57 in54 sn57 11140.846016
Rwneg54_58 in54 sn58 3183.098862
Rwneg54_59 in54 sn59 11140.846016
Rwneg54_60 in54 sn60 11140.846016
Rwneg54_61 in54 sn61 3183.098862
Rwneg54_62 in54 sn62 11140.846016
Rwneg54_63 in54 sn63 3183.098862
Rwneg54_64 in54 sn64 3183.098862
Rwneg54_65 in54 sn65 3183.098862
Rwneg54_66 in54 sn66 3183.098862
Rwneg54_67 in54 sn67 3183.098862
Rwneg54_68 in54 sn68 11140.846016
Rwneg54_69 in54 sn69 3183.098862
Rwneg54_70 in54 sn70 3183.098862
Rwneg54_71 in54 sn71 11140.846016
Rwneg54_72 in54 sn72 11140.846016
Rwneg54_73 in54 sn73 11140.846016
Rwneg54_74 in54 sn74 11140.846016
Rwneg54_75 in54 sn75 3183.098862
Rwneg54_76 in54 sn76 3183.098862
Rwneg54_77 in54 sn77 3183.098862
Rwneg54_78 in54 sn78 3183.098862
Rwneg54_79 in54 sn79 11140.846016
Rwneg54_80 in54 sn80 3183.098862
Rwneg54_81 in54 sn81 3183.098862
Rwneg54_82 in54 sn82 11140.846016
Rwneg54_83 in54 sn83 3183.098862
Rwneg54_84 in54 sn84 11140.846016
Rwneg54_85 in54 sn85 11140.846016
Rwneg54_86 in54 sn86 11140.846016
Rwneg54_87 in54 sn87 3183.098862
Rwneg54_88 in54 sn88 3183.098862
Rwneg54_89 in54 sn89 3183.098862
Rwneg54_90 in54 sn90 3183.098862
Rwneg54_91 in54 sn91 11140.846016
Rwneg54_92 in54 sn92 11140.846016
Rwneg54_93 in54 sn93 3183.098862
Rwneg54_94 in54 sn94 11140.846016
Rwneg54_95 in54 sn95 3183.098862
Rwneg54_96 in54 sn96 3183.098862
Rwneg54_97 in54 sn97 11140.846016
Rwneg54_98 in54 sn98 11140.846016
Rwneg54_99 in54 sn99 3183.098862
Rwneg54_100 in54 sn100 3183.098862
Rwneg55_1 in55 sn1 3183.098862
Rwneg55_2 in55 sn2 11140.846016
Rwneg55_3 in55 sn3 3183.098862
Rwneg55_4 in55 sn4 3183.098862
Rwneg55_5 in55 sn5 11140.846016
Rwneg55_6 in55 sn6 3183.098862
Rwneg55_7 in55 sn7 3183.098862
Rwneg55_8 in55 sn8 11140.846016
Rwneg55_9 in55 sn9 11140.846016
Rwneg55_10 in55 sn10 3183.098862
Rwneg55_11 in55 sn11 3183.098862
Rwneg55_12 in55 sn12 3183.098862
Rwneg55_13 in55 sn13 11140.846016
Rwneg55_14 in55 sn14 11140.846016
Rwneg55_15 in55 sn15 3183.098862
Rwneg55_16 in55 sn16 3183.098862
Rwneg55_17 in55 sn17 3183.098862
Rwneg55_18 in55 sn18 3183.098862
Rwneg55_19 in55 sn19 3183.098862
Rwneg55_20 in55 sn20 11140.846016
Rwneg55_21 in55 sn21 3183.098862
Rwneg55_22 in55 sn22 11140.846016
Rwneg55_23 in55 sn23 3183.098862
Rwneg55_24 in55 sn24 11140.846016
Rwneg55_25 in55 sn25 3183.098862
Rwneg55_26 in55 sn26 3183.098862
Rwneg55_27 in55 sn27 11140.846016
Rwneg55_28 in55 sn28 11140.846016
Rwneg55_29 in55 sn29 11140.846016
Rwneg55_30 in55 sn30 3183.098862
Rwneg55_31 in55 sn31 11140.846016
Rwneg55_32 in55 sn32 3183.098862
Rwneg55_33 in55 sn33 3183.098862
Rwneg55_34 in55 sn34 3183.098862
Rwneg55_35 in55 sn35 11140.846016
Rwneg55_36 in55 sn36 3183.098862
Rwneg55_37 in55 sn37 3183.098862
Rwneg55_38 in55 sn38 11140.846016
Rwneg55_39 in55 sn39 11140.846016
Rwneg55_40 in55 sn40 3183.098862
Rwneg55_41 in55 sn41 3183.098862
Rwneg55_42 in55 sn42 3183.098862
Rwneg55_43 in55 sn43 11140.846016
Rwneg55_44 in55 sn44 3183.098862
Rwneg55_45 in55 sn45 3183.098862
Rwneg55_46 in55 sn46 3183.098862
Rwneg55_47 in55 sn47 11140.846016
Rwneg55_48 in55 sn48 3183.098862
Rwneg55_49 in55 sn49 11140.846016
Rwneg55_50 in55 sn50 11140.846016
Rwneg55_51 in55 sn51 3183.098862
Rwneg55_52 in55 sn52 3183.098862
Rwneg55_53 in55 sn53 3183.098862
Rwneg55_54 in55 sn54 11140.846016
Rwneg55_55 in55 sn55 11140.846016
Rwneg55_56 in55 sn56 3183.098862
Rwneg55_57 in55 sn57 3183.098862
Rwneg55_58 in55 sn58 11140.846016
Rwneg55_59 in55 sn59 3183.098862
Rwneg55_60 in55 sn60 3183.098862
Rwneg55_61 in55 sn61 3183.098862
Rwneg55_62 in55 sn62 3183.098862
Rwneg55_63 in55 sn63 3183.098862
Rwneg55_64 in55 sn64 3183.098862
Rwneg55_65 in55 sn65 11140.846016
Rwneg55_66 in55 sn66 3183.098862
Rwneg55_67 in55 sn67 11140.846016
Rwneg55_68 in55 sn68 11140.846016
Rwneg55_69 in55 sn69 3183.098862
Rwneg55_70 in55 sn70 11140.846016
Rwneg55_71 in55 sn71 3183.098862
Rwneg55_72 in55 sn72 11140.846016
Rwneg55_73 in55 sn73 11140.846016
Rwneg55_74 in55 sn74 3183.098862
Rwneg55_75 in55 sn75 3183.098862
Rwneg55_76 in55 sn76 3183.098862
Rwneg55_77 in55 sn77 11140.846016
Rwneg55_78 in55 sn78 3183.098862
Rwneg55_79 in55 sn79 3183.098862
Rwneg55_80 in55 sn80 3183.098862
Rwneg55_81 in55 sn81 3183.098862
Rwneg55_82 in55 sn82 3183.098862
Rwneg55_83 in55 sn83 11140.846016
Rwneg55_84 in55 sn84 11140.846016
Rwneg55_85 in55 sn85 3183.098862
Rwneg55_86 in55 sn86 3183.098862
Rwneg55_87 in55 sn87 11140.846016
Rwneg55_88 in55 sn88 11140.846016
Rwneg55_89 in55 sn89 11140.846016
Rwneg55_90 in55 sn90 11140.846016
Rwneg55_91 in55 sn91 3183.098862
Rwneg55_92 in55 sn92 11140.846016
Rwneg55_93 in55 sn93 3183.098862
Rwneg55_94 in55 sn94 11140.846016
Rwneg55_95 in55 sn95 11140.846016
Rwneg55_96 in55 sn96 3183.098862
Rwneg55_97 in55 sn97 3183.098862
Rwneg55_98 in55 sn98 11140.846016
Rwneg55_99 in55 sn99 11140.846016
Rwneg55_100 in55 sn100 11140.846016
Rwneg56_1 in56 sn1 3183.098862
Rwneg56_2 in56 sn2 11140.846016
Rwneg56_3 in56 sn3 11140.846016
Rwneg56_4 in56 sn4 11140.846016
Rwneg56_5 in56 sn5 11140.846016
Rwneg56_6 in56 sn6 3183.098862
Rwneg56_7 in56 sn7 3183.098862
Rwneg56_8 in56 sn8 11140.846016
Rwneg56_9 in56 sn9 3183.098862
Rwneg56_10 in56 sn10 3183.098862
Rwneg56_11 in56 sn11 3183.098862
Rwneg56_12 in56 sn12 3183.098862
Rwneg56_13 in56 sn13 3183.098862
Rwneg56_14 in56 sn14 3183.098862
Rwneg56_15 in56 sn15 11140.846016
Rwneg56_16 in56 sn16 11140.846016
Rwneg56_17 in56 sn17 3183.098862
Rwneg56_18 in56 sn18 11140.846016
Rwneg56_19 in56 sn19 3183.098862
Rwneg56_20 in56 sn20 11140.846016
Rwneg56_21 in56 sn21 11140.846016
Rwneg56_22 in56 sn22 11140.846016
Rwneg56_23 in56 sn23 3183.098862
Rwneg56_24 in56 sn24 11140.846016
Rwneg56_25 in56 sn25 11140.846016
Rwneg56_26 in56 sn26 11140.846016
Rwneg56_27 in56 sn27 3183.098862
Rwneg56_28 in56 sn28 3183.098862
Rwneg56_29 in56 sn29 3183.098862
Rwneg56_30 in56 sn30 3183.098862
Rwneg56_31 in56 sn31 11140.846016
Rwneg56_32 in56 sn32 11140.846016
Rwneg56_33 in56 sn33 3183.098862
Rwneg56_34 in56 sn34 11140.846016
Rwneg56_35 in56 sn35 3183.098862
Rwneg56_36 in56 sn36 11140.846016
Rwneg56_37 in56 sn37 11140.846016
Rwneg56_38 in56 sn38 11140.846016
Rwneg56_39 in56 sn39 11140.846016
Rwneg56_40 in56 sn40 11140.846016
Rwneg56_41 in56 sn41 11140.846016
Rwneg56_42 in56 sn42 3183.098862
Rwneg56_43 in56 sn43 11140.846016
Rwneg56_44 in56 sn44 3183.098862
Rwneg56_45 in56 sn45 3183.098862
Rwneg56_46 in56 sn46 3183.098862
Rwneg56_47 in56 sn47 11140.846016
Rwneg56_48 in56 sn48 11140.846016
Rwneg56_49 in56 sn49 3183.098862
Rwneg56_50 in56 sn50 3183.098862
Rwneg56_51 in56 sn51 11140.846016
Rwneg56_52 in56 sn52 11140.846016
Rwneg56_53 in56 sn53 11140.846016
Rwneg56_54 in56 sn54 3183.098862
Rwneg56_55 in56 sn55 3183.098862
Rwneg56_56 in56 sn56 11140.846016
Rwneg56_57 in56 sn57 3183.098862
Rwneg56_58 in56 sn58 3183.098862
Rwneg56_59 in56 sn59 11140.846016
Rwneg56_60 in56 sn60 3183.098862
Rwneg56_61 in56 sn61 3183.098862
Rwneg56_62 in56 sn62 3183.098862
Rwneg56_63 in56 sn63 11140.846016
Rwneg56_64 in56 sn64 11140.846016
Rwneg56_65 in56 sn65 3183.098862
Rwneg56_66 in56 sn66 11140.846016
Rwneg56_67 in56 sn67 11140.846016
Rwneg56_68 in56 sn68 11140.846016
Rwneg56_69 in56 sn69 11140.846016
Rwneg56_70 in56 sn70 3183.098862
Rwneg56_71 in56 sn71 11140.846016
Rwneg56_72 in56 sn72 11140.846016
Rwneg56_73 in56 sn73 11140.846016
Rwneg56_74 in56 sn74 3183.098862
Rwneg56_75 in56 sn75 11140.846016
Rwneg56_76 in56 sn76 3183.098862
Rwneg56_77 in56 sn77 3183.098862
Rwneg56_78 in56 sn78 3183.098862
Rwneg56_79 in56 sn79 11140.846016
Rwneg56_80 in56 sn80 11140.846016
Rwneg56_81 in56 sn81 3183.098862
Rwneg56_82 in56 sn82 11140.846016
Rwneg56_83 in56 sn83 11140.846016
Rwneg56_84 in56 sn84 11140.846016
Rwneg56_85 in56 sn85 3183.098862
Rwneg56_86 in56 sn86 3183.098862
Rwneg56_87 in56 sn87 3183.098862
Rwneg56_88 in56 sn88 11140.846016
Rwneg56_89 in56 sn89 11140.846016
Rwneg56_90 in56 sn90 3183.098862
Rwneg56_91 in56 sn91 3183.098862
Rwneg56_92 in56 sn92 11140.846016
Rwneg56_93 in56 sn93 3183.098862
Rwneg56_94 in56 sn94 3183.098862
Rwneg56_95 in56 sn95 11140.846016
Rwneg56_96 in56 sn96 11140.846016
Rwneg56_97 in56 sn97 3183.098862
Rwneg56_98 in56 sn98 3183.098862
Rwneg56_99 in56 sn99 11140.846016
Rwneg56_100 in56 sn100 11140.846016
Rwneg57_1 in57 sn1 11140.846016
Rwneg57_2 in57 sn2 3183.098862
Rwneg57_3 in57 sn3 3183.098862
Rwneg57_4 in57 sn4 3183.098862
Rwneg57_5 in57 sn5 11140.846016
Rwneg57_6 in57 sn6 3183.098862
Rwneg57_7 in57 sn7 3183.098862
Rwneg57_8 in57 sn8 11140.846016
Rwneg57_9 in57 sn9 11140.846016
Rwneg57_10 in57 sn10 11140.846016
Rwneg57_11 in57 sn11 11140.846016
Rwneg57_12 in57 sn12 11140.846016
Rwneg57_13 in57 sn13 3183.098862
Rwneg57_14 in57 sn14 3183.098862
Rwneg57_15 in57 sn15 11140.846016
Rwneg57_16 in57 sn16 11140.846016
Rwneg57_17 in57 sn17 3183.098862
Rwneg57_18 in57 sn18 3183.098862
Rwneg57_19 in57 sn19 3183.098862
Rwneg57_20 in57 sn20 3183.098862
Rwneg57_21 in57 sn21 11140.846016
Rwneg57_22 in57 sn22 3183.098862
Rwneg57_23 in57 sn23 3183.098862
Rwneg57_24 in57 sn24 3183.098862
Rwneg57_25 in57 sn25 11140.846016
Rwneg57_26 in57 sn26 11140.846016
Rwneg57_27 in57 sn27 11140.846016
Rwneg57_28 in57 sn28 11140.846016
Rwneg57_29 in57 sn29 11140.846016
Rwneg57_30 in57 sn30 3183.098862
Rwneg57_31 in57 sn31 11140.846016
Rwneg57_32 in57 sn32 11140.846016
Rwneg57_33 in57 sn33 3183.098862
Rwneg57_34 in57 sn34 3183.098862
Rwneg57_35 in57 sn35 3183.098862
Rwneg57_36 in57 sn36 11140.846016
Rwneg57_37 in57 sn37 11140.846016
Rwneg57_38 in57 sn38 3183.098862
Rwneg57_39 in57 sn39 11140.846016
Rwneg57_40 in57 sn40 3183.098862
Rwneg57_41 in57 sn41 11140.846016
Rwneg57_42 in57 sn42 3183.098862
Rwneg57_43 in57 sn43 3183.098862
Rwneg57_44 in57 sn44 11140.846016
Rwneg57_45 in57 sn45 11140.846016
Rwneg57_46 in57 sn46 3183.098862
Rwneg57_47 in57 sn47 11140.846016
Rwneg57_48 in57 sn48 11140.846016
Rwneg57_49 in57 sn49 3183.098862
Rwneg57_50 in57 sn50 3183.098862
Rwneg57_51 in57 sn51 11140.846016
Rwneg57_52 in57 sn52 3183.098862
Rwneg57_53 in57 sn53 3183.098862
Rwneg57_54 in57 sn54 3183.098862
Rwneg57_55 in57 sn55 11140.846016
Rwneg57_56 in57 sn56 3183.098862
Rwneg57_57 in57 sn57 11140.846016
Rwneg57_58 in57 sn58 11140.846016
Rwneg57_59 in57 sn59 3183.098862
Rwneg57_60 in57 sn60 11140.846016
Rwneg57_61 in57 sn61 11140.846016
Rwneg57_62 in57 sn62 11140.846016
Rwneg57_63 in57 sn63 3183.098862
Rwneg57_64 in57 sn64 11140.846016
Rwneg57_65 in57 sn65 11140.846016
Rwneg57_66 in57 sn66 11140.846016
Rwneg57_67 in57 sn67 3183.098862
Rwneg57_68 in57 sn68 3183.098862
Rwneg57_69 in57 sn69 3183.098862
Rwneg57_70 in57 sn70 3183.098862
Rwneg57_71 in57 sn71 11140.846016
Rwneg57_72 in57 sn72 3183.098862
Rwneg57_73 in57 sn73 11140.846016
Rwneg57_74 in57 sn74 11140.846016
Rwneg57_75 in57 sn75 11140.846016
Rwneg57_76 in57 sn76 11140.846016
Rwneg57_77 in57 sn77 3183.098862
Rwneg57_78 in57 sn78 3183.098862
Rwneg57_79 in57 sn79 11140.846016
Rwneg57_80 in57 sn80 11140.846016
Rwneg57_81 in57 sn81 11140.846016
Rwneg57_82 in57 sn82 11140.846016
Rwneg57_83 in57 sn83 3183.098862
Rwneg57_84 in57 sn84 11140.846016
Rwneg57_85 in57 sn85 11140.846016
Rwneg57_86 in57 sn86 11140.846016
Rwneg57_87 in57 sn87 11140.846016
Rwneg57_88 in57 sn88 11140.846016
Rwneg57_89 in57 sn89 11140.846016
Rwneg57_90 in57 sn90 3183.098862
Rwneg57_91 in57 sn91 3183.098862
Rwneg57_92 in57 sn92 3183.098862
Rwneg57_93 in57 sn93 3183.098862
Rwneg57_94 in57 sn94 3183.098862
Rwneg57_95 in57 sn95 11140.846016
Rwneg57_96 in57 sn96 3183.098862
Rwneg57_97 in57 sn97 11140.846016
Rwneg57_98 in57 sn98 11140.846016
Rwneg57_99 in57 sn99 3183.098862
Rwneg57_100 in57 sn100 3183.098862
Rwneg58_1 in58 sn1 11140.846016
Rwneg58_2 in58 sn2 3183.098862
Rwneg58_3 in58 sn3 11140.846016
Rwneg58_4 in58 sn4 11140.846016
Rwneg58_5 in58 sn5 11140.846016
Rwneg58_6 in58 sn6 11140.846016
Rwneg58_7 in58 sn7 11140.846016
Rwneg58_8 in58 sn8 11140.846016
Rwneg58_9 in58 sn9 11140.846016
Rwneg58_10 in58 sn10 3183.098862
Rwneg58_11 in58 sn11 3183.098862
Rwneg58_12 in58 sn12 3183.098862
Rwneg58_13 in58 sn13 11140.846016
Rwneg58_14 in58 sn14 11140.846016
Rwneg58_15 in58 sn15 3183.098862
Rwneg58_16 in58 sn16 3183.098862
Rwneg58_17 in58 sn17 3183.098862
Rwneg58_18 in58 sn18 11140.846016
Rwneg58_19 in58 sn19 11140.846016
Rwneg58_20 in58 sn20 3183.098862
Rwneg58_21 in58 sn21 11140.846016
Rwneg58_22 in58 sn22 11140.846016
Rwneg58_23 in58 sn23 11140.846016
Rwneg58_24 in58 sn24 11140.846016
Rwneg58_25 in58 sn25 11140.846016
Rwneg58_26 in58 sn26 3183.098862
Rwneg58_27 in58 sn27 3183.098862
Rwneg58_28 in58 sn28 3183.098862
Rwneg58_29 in58 sn29 11140.846016
Rwneg58_30 in58 sn30 11140.846016
Rwneg58_31 in58 sn31 3183.098862
Rwneg58_32 in58 sn32 3183.098862
Rwneg58_33 in58 sn33 11140.846016
Rwneg58_34 in58 sn34 3183.098862
Rwneg58_35 in58 sn35 11140.846016
Rwneg58_36 in58 sn36 11140.846016
Rwneg58_37 in58 sn37 11140.846016
Rwneg58_38 in58 sn38 3183.098862
Rwneg58_39 in58 sn39 11140.846016
Rwneg58_40 in58 sn40 3183.098862
Rwneg58_41 in58 sn41 11140.846016
Rwneg58_42 in58 sn42 3183.098862
Rwneg58_43 in58 sn43 3183.098862
Rwneg58_44 in58 sn44 11140.846016
Rwneg58_45 in58 sn45 11140.846016
Rwneg58_46 in58 sn46 11140.846016
Rwneg58_47 in58 sn47 3183.098862
Rwneg58_48 in58 sn48 11140.846016
Rwneg58_49 in58 sn49 11140.846016
Rwneg58_50 in58 sn50 3183.098862
Rwneg58_51 in58 sn51 11140.846016
Rwneg58_52 in58 sn52 11140.846016
Rwneg58_53 in58 sn53 3183.098862
Rwneg58_54 in58 sn54 3183.098862
Rwneg58_55 in58 sn55 11140.846016
Rwneg58_56 in58 sn56 3183.098862
Rwneg58_57 in58 sn57 11140.846016
Rwneg58_58 in58 sn58 11140.846016
Rwneg58_59 in58 sn59 3183.098862
Rwneg58_60 in58 sn60 11140.846016
Rwneg58_61 in58 sn61 3183.098862
Rwneg58_62 in58 sn62 3183.098862
Rwneg58_63 in58 sn63 3183.098862
Rwneg58_64 in58 sn64 3183.098862
Rwneg58_65 in58 sn65 11140.846016
Rwneg58_66 in58 sn66 11140.846016
Rwneg58_67 in58 sn67 11140.846016
Rwneg58_68 in58 sn68 3183.098862
Rwneg58_69 in58 sn69 3183.098862
Rwneg58_70 in58 sn70 3183.098862
Rwneg58_71 in58 sn71 3183.098862
Rwneg58_72 in58 sn72 3183.098862
Rwneg58_73 in58 sn73 11140.846016
Rwneg58_74 in58 sn74 11140.846016
Rwneg58_75 in58 sn75 3183.098862
Rwneg58_76 in58 sn76 11140.846016
Rwneg58_77 in58 sn77 11140.846016
Rwneg58_78 in58 sn78 11140.846016
Rwneg58_79 in58 sn79 11140.846016
Rwneg58_80 in58 sn80 11140.846016
Rwneg58_81 in58 sn81 3183.098862
Rwneg58_82 in58 sn82 3183.098862
Rwneg58_83 in58 sn83 11140.846016
Rwneg58_84 in58 sn84 11140.846016
Rwneg58_85 in58 sn85 3183.098862
Rwneg58_86 in58 sn86 3183.098862
Rwneg58_87 in58 sn87 11140.846016
Rwneg58_88 in58 sn88 11140.846016
Rwneg58_89 in58 sn89 11140.846016
Rwneg58_90 in58 sn90 3183.098862
Rwneg58_91 in58 sn91 11140.846016
Rwneg58_92 in58 sn92 11140.846016
Rwneg58_93 in58 sn93 11140.846016
Rwneg58_94 in58 sn94 11140.846016
Rwneg58_95 in58 sn95 11140.846016
Rwneg58_96 in58 sn96 3183.098862
Rwneg58_97 in58 sn97 11140.846016
Rwneg58_98 in58 sn98 3183.098862
Rwneg58_99 in58 sn99 11140.846016
Rwneg58_100 in58 sn100 11140.846016
Rwneg59_1 in59 sn1 11140.846016
Rwneg59_2 in59 sn2 11140.846016
Rwneg59_3 in59 sn3 11140.846016
Rwneg59_4 in59 sn4 3183.098862
Rwneg59_5 in59 sn5 11140.846016
Rwneg59_6 in59 sn6 11140.846016
Rwneg59_7 in59 sn7 3183.098862
Rwneg59_8 in59 sn8 11140.846016
Rwneg59_9 in59 sn9 3183.098862
Rwneg59_10 in59 sn10 11140.846016
Rwneg59_11 in59 sn11 11140.846016
Rwneg59_12 in59 sn12 11140.846016
Rwneg59_13 in59 sn13 3183.098862
Rwneg59_14 in59 sn14 11140.846016
Rwneg59_15 in59 sn15 3183.098862
Rwneg59_16 in59 sn16 11140.846016
Rwneg59_17 in59 sn17 3183.098862
Rwneg59_18 in59 sn18 11140.846016
Rwneg59_19 in59 sn19 3183.098862
Rwneg59_20 in59 sn20 11140.846016
Rwneg59_21 in59 sn21 3183.098862
Rwneg59_22 in59 sn22 3183.098862
Rwneg59_23 in59 sn23 11140.846016
Rwneg59_24 in59 sn24 11140.846016
Rwneg59_25 in59 sn25 11140.846016
Rwneg59_26 in59 sn26 3183.098862
Rwneg59_27 in59 sn27 3183.098862
Rwneg59_28 in59 sn28 11140.846016
Rwneg59_29 in59 sn29 3183.098862
Rwneg59_30 in59 sn30 11140.846016
Rwneg59_31 in59 sn31 11140.846016
Rwneg59_32 in59 sn32 11140.846016
Rwneg59_33 in59 sn33 11140.846016
Rwneg59_34 in59 sn34 11140.846016
Rwneg59_35 in59 sn35 3183.098862
Rwneg59_36 in59 sn36 11140.846016
Rwneg59_37 in59 sn37 11140.846016
Rwneg59_38 in59 sn38 11140.846016
Rwneg59_39 in59 sn39 11140.846016
Rwneg59_40 in59 sn40 11140.846016
Rwneg59_41 in59 sn41 11140.846016
Rwneg59_42 in59 sn42 3183.098862
Rwneg59_43 in59 sn43 3183.098862
Rwneg59_44 in59 sn44 11140.846016
Rwneg59_45 in59 sn45 3183.098862
Rwneg59_46 in59 sn46 3183.098862
Rwneg59_47 in59 sn47 3183.098862
Rwneg59_48 in59 sn48 11140.846016
Rwneg59_49 in59 sn49 11140.846016
Rwneg59_50 in59 sn50 11140.846016
Rwneg59_51 in59 sn51 3183.098862
Rwneg59_52 in59 sn52 3183.098862
Rwneg59_53 in59 sn53 11140.846016
Rwneg59_54 in59 sn54 11140.846016
Rwneg59_55 in59 sn55 3183.098862
Rwneg59_56 in59 sn56 11140.846016
Rwneg59_57 in59 sn57 11140.846016
Rwneg59_58 in59 sn58 3183.098862
Rwneg59_59 in59 sn59 3183.098862
Rwneg59_60 in59 sn60 11140.846016
Rwneg59_61 in59 sn61 11140.846016
Rwneg59_62 in59 sn62 11140.846016
Rwneg59_63 in59 sn63 11140.846016
Rwneg59_64 in59 sn64 11140.846016
Rwneg59_65 in59 sn65 11140.846016
Rwneg59_66 in59 sn66 11140.846016
Rwneg59_67 in59 sn67 3183.098862
Rwneg59_68 in59 sn68 3183.098862
Rwneg59_69 in59 sn69 11140.846016
Rwneg59_70 in59 sn70 3183.098862
Rwneg59_71 in59 sn71 11140.846016
Rwneg59_72 in59 sn72 11140.846016
Rwneg59_73 in59 sn73 11140.846016
Rwneg59_74 in59 sn74 11140.846016
Rwneg59_75 in59 sn75 3183.098862
Rwneg59_76 in59 sn76 3183.098862
Rwneg59_77 in59 sn77 3183.098862
Rwneg59_78 in59 sn78 3183.098862
Rwneg59_79 in59 sn79 11140.846016
Rwneg59_80 in59 sn80 11140.846016
Rwneg59_81 in59 sn81 11140.846016
Rwneg59_82 in59 sn82 3183.098862
Rwneg59_83 in59 sn83 11140.846016
Rwneg59_84 in59 sn84 11140.846016
Rwneg59_85 in59 sn85 3183.098862
Rwneg59_86 in59 sn86 11140.846016
Rwneg59_87 in59 sn87 11140.846016
Rwneg59_88 in59 sn88 11140.846016
Rwneg59_89 in59 sn89 11140.846016
Rwneg59_90 in59 sn90 3183.098862
Rwneg59_91 in59 sn91 3183.098862
Rwneg59_92 in59 sn92 11140.846016
Rwneg59_93 in59 sn93 11140.846016
Rwneg59_94 in59 sn94 11140.846016
Rwneg59_95 in59 sn95 3183.098862
Rwneg59_96 in59 sn96 3183.098862
Rwneg59_97 in59 sn97 3183.098862
Rwneg59_98 in59 sn98 11140.846016
Rwneg59_99 in59 sn99 11140.846016
Rwneg59_100 in59 sn100 11140.846016
Rwneg60_1 in60 sn1 3183.098862
Rwneg60_2 in60 sn2 11140.846016
Rwneg60_3 in60 sn3 3183.098862
Rwneg60_4 in60 sn4 11140.846016
Rwneg60_5 in60 sn5 3183.098862
Rwneg60_6 in60 sn6 11140.846016
Rwneg60_7 in60 sn7 3183.098862
Rwneg60_8 in60 sn8 3183.098862
Rwneg60_9 in60 sn9 11140.846016
Rwneg60_10 in60 sn10 3183.098862
Rwneg60_11 in60 sn11 3183.098862
Rwneg60_12 in60 sn12 3183.098862
Rwneg60_13 in60 sn13 3183.098862
Rwneg60_14 in60 sn14 3183.098862
Rwneg60_15 in60 sn15 11140.846016
Rwneg60_16 in60 sn16 3183.098862
Rwneg60_17 in60 sn17 11140.846016
Rwneg60_18 in60 sn18 11140.846016
Rwneg60_19 in60 sn19 11140.846016
Rwneg60_20 in60 sn20 11140.846016
Rwneg60_21 in60 sn21 11140.846016
Rwneg60_22 in60 sn22 11140.846016
Rwneg60_23 in60 sn23 3183.098862
Rwneg60_24 in60 sn24 3183.098862
Rwneg60_25 in60 sn25 11140.846016
Rwneg60_26 in60 sn26 3183.098862
Rwneg60_27 in60 sn27 11140.846016
Rwneg60_28 in60 sn28 3183.098862
Rwneg60_29 in60 sn29 11140.846016
Rwneg60_30 in60 sn30 3183.098862
Rwneg60_31 in60 sn31 11140.846016
Rwneg60_32 in60 sn32 11140.846016
Rwneg60_33 in60 sn33 11140.846016
Rwneg60_34 in60 sn34 11140.846016
Rwneg60_35 in60 sn35 3183.098862
Rwneg60_36 in60 sn36 11140.846016
Rwneg60_37 in60 sn37 11140.846016
Rwneg60_38 in60 sn38 11140.846016
Rwneg60_39 in60 sn39 3183.098862
Rwneg60_40 in60 sn40 3183.098862
Rwneg60_41 in60 sn41 11140.846016
Rwneg60_42 in60 sn42 3183.098862
Rwneg60_43 in60 sn43 11140.846016
Rwneg60_44 in60 sn44 3183.098862
Rwneg60_45 in60 sn45 3183.098862
Rwneg60_46 in60 sn46 3183.098862
Rwneg60_47 in60 sn47 11140.846016
Rwneg60_48 in60 sn48 11140.846016
Rwneg60_49 in60 sn49 11140.846016
Rwneg60_50 in60 sn50 11140.846016
Rwneg60_51 in60 sn51 11140.846016
Rwneg60_52 in60 sn52 11140.846016
Rwneg60_53 in60 sn53 11140.846016
Rwneg60_54 in60 sn54 3183.098862
Rwneg60_55 in60 sn55 3183.098862
Rwneg60_56 in60 sn56 3183.098862
Rwneg60_57 in60 sn57 11140.846016
Rwneg60_58 in60 sn58 3183.098862
Rwneg60_59 in60 sn59 11140.846016
Rwneg60_60 in60 sn60 3183.098862
Rwneg60_61 in60 sn61 11140.846016
Rwneg60_62 in60 sn62 3183.098862
Rwneg60_63 in60 sn63 11140.846016
Rwneg60_64 in60 sn64 11140.846016
Rwneg60_65 in60 sn65 11140.846016
Rwneg60_66 in60 sn66 11140.846016
Rwneg60_67 in60 sn67 11140.846016
Rwneg60_68 in60 sn68 11140.846016
Rwneg60_69 in60 sn69 11140.846016
Rwneg60_70 in60 sn70 3183.098862
Rwneg60_71 in60 sn71 3183.098862
Rwneg60_72 in60 sn72 11140.846016
Rwneg60_73 in60 sn73 11140.846016
Rwneg60_74 in60 sn74 11140.846016
Rwneg60_75 in60 sn75 3183.098862
Rwneg60_76 in60 sn76 3183.098862
Rwneg60_77 in60 sn77 3183.098862
Rwneg60_78 in60 sn78 3183.098862
Rwneg60_79 in60 sn79 11140.846016
Rwneg60_80 in60 sn80 11140.846016
Rwneg60_81 in60 sn81 3183.098862
Rwneg60_82 in60 sn82 11140.846016
Rwneg60_83 in60 sn83 11140.846016
Rwneg60_84 in60 sn84 11140.846016
Rwneg60_85 in60 sn85 11140.846016
Rwneg60_86 in60 sn86 3183.098862
Rwneg60_87 in60 sn87 3183.098862
Rwneg60_88 in60 sn88 11140.846016
Rwneg60_89 in60 sn89 11140.846016
Rwneg60_90 in60 sn90 3183.098862
Rwneg60_91 in60 sn91 3183.098862
Rwneg60_92 in60 sn92 3183.098862
Rwneg60_93 in60 sn93 3183.098862
Rwneg60_94 in60 sn94 3183.098862
Rwneg60_95 in60 sn95 11140.846016
Rwneg60_96 in60 sn96 11140.846016
Rwneg60_97 in60 sn97 11140.846016
Rwneg60_98 in60 sn98 11140.846016
Rwneg60_99 in60 sn99 3183.098862
Rwneg60_100 in60 sn100 11140.846016
Rwneg61_1 in61 sn1 11140.846016
Rwneg61_2 in61 sn2 3183.098862
Rwneg61_3 in61 sn3 11140.846016
Rwneg61_4 in61 sn4 11140.846016
Rwneg61_5 in61 sn5 11140.846016
Rwneg61_6 in61 sn6 3183.098862
Rwneg61_7 in61 sn7 3183.098862
Rwneg61_8 in61 sn8 3183.098862
Rwneg61_9 in61 sn9 3183.098862
Rwneg61_10 in61 sn10 3183.098862
Rwneg61_11 in61 sn11 11140.846016
Rwneg61_12 in61 sn12 11140.846016
Rwneg61_13 in61 sn13 3183.098862
Rwneg61_14 in61 sn14 11140.846016
Rwneg61_15 in61 sn15 11140.846016
Rwneg61_16 in61 sn16 11140.846016
Rwneg61_17 in61 sn17 11140.846016
Rwneg61_18 in61 sn18 3183.098862
Rwneg61_19 in61 sn19 3183.098862
Rwneg61_20 in61 sn20 11140.846016
Rwneg61_21 in61 sn21 11140.846016
Rwneg61_22 in61 sn22 3183.098862
Rwneg61_23 in61 sn23 11140.846016
Rwneg61_24 in61 sn24 11140.846016
Rwneg61_25 in61 sn25 3183.098862
Rwneg61_26 in61 sn26 3183.098862
Rwneg61_27 in61 sn27 3183.098862
Rwneg61_28 in61 sn28 11140.846016
Rwneg61_29 in61 sn29 3183.098862
Rwneg61_30 in61 sn30 11140.846016
Rwneg61_31 in61 sn31 11140.846016
Rwneg61_32 in61 sn32 11140.846016
Rwneg61_33 in61 sn33 3183.098862
Rwneg61_34 in61 sn34 3183.098862
Rwneg61_35 in61 sn35 3183.098862
Rwneg61_36 in61 sn36 11140.846016
Rwneg61_37 in61 sn37 11140.846016
Rwneg61_38 in61 sn38 3183.098862
Rwneg61_39 in61 sn39 3183.098862
Rwneg61_40 in61 sn40 11140.846016
Rwneg61_41 in61 sn41 11140.846016
Rwneg61_42 in61 sn42 3183.098862
Rwneg61_43 in61 sn43 3183.098862
Rwneg61_44 in61 sn44 11140.846016
Rwneg61_45 in61 sn45 3183.098862
Rwneg61_46 in61 sn46 3183.098862
Rwneg61_47 in61 sn47 11140.846016
Rwneg61_48 in61 sn48 11140.846016
Rwneg61_49 in61 sn49 11140.846016
Rwneg61_50 in61 sn50 11140.846016
Rwneg61_51 in61 sn51 3183.098862
Rwneg61_52 in61 sn52 3183.098862
Rwneg61_53 in61 sn53 11140.846016
Rwneg61_54 in61 sn54 3183.098862
Rwneg61_55 in61 sn55 3183.098862
Rwneg61_56 in61 sn56 3183.098862
Rwneg61_57 in61 sn57 11140.846016
Rwneg61_58 in61 sn58 11140.846016
Rwneg61_59 in61 sn59 11140.846016
Rwneg61_60 in61 sn60 11140.846016
Rwneg61_61 in61 sn61 3183.098862
Rwneg61_62 in61 sn62 3183.098862
Rwneg61_63 in61 sn63 11140.846016
Rwneg61_64 in61 sn64 11140.846016
Rwneg61_65 in61 sn65 11140.846016
Rwneg61_66 in61 sn66 3183.098862
Rwneg61_67 in61 sn67 3183.098862
Rwneg61_68 in61 sn68 11140.846016
Rwneg61_69 in61 sn69 11140.846016
Rwneg61_70 in61 sn70 3183.098862
Rwneg61_71 in61 sn71 3183.098862
Rwneg61_72 in61 sn72 3183.098862
Rwneg61_73 in61 sn73 11140.846016
Rwneg61_74 in61 sn74 11140.846016
Rwneg61_75 in61 sn75 11140.846016
Rwneg61_76 in61 sn76 11140.846016
Rwneg61_77 in61 sn77 11140.846016
Rwneg61_78 in61 sn78 3183.098862
Rwneg61_79 in61 sn79 11140.846016
Rwneg61_80 in61 sn80 11140.846016
Rwneg61_81 in61 sn81 3183.098862
Rwneg61_82 in61 sn82 11140.846016
Rwneg61_83 in61 sn83 3183.098862
Rwneg61_84 in61 sn84 11140.846016
Rwneg61_85 in61 sn85 11140.846016
Rwneg61_86 in61 sn86 3183.098862
Rwneg61_87 in61 sn87 11140.846016
Rwneg61_88 in61 sn88 3183.098862
Rwneg61_89 in61 sn89 11140.846016
Rwneg61_90 in61 sn90 3183.098862
Rwneg61_91 in61 sn91 11140.846016
Rwneg61_92 in61 sn92 11140.846016
Rwneg61_93 in61 sn93 3183.098862
Rwneg61_94 in61 sn94 11140.846016
Rwneg61_95 in61 sn95 11140.846016
Rwneg61_96 in61 sn96 11140.846016
Rwneg61_97 in61 sn97 11140.846016
Rwneg61_98 in61 sn98 11140.846016
Rwneg61_99 in61 sn99 3183.098862
Rwneg61_100 in61 sn100 11140.846016
Rwneg62_1 in62 sn1 3183.098862
Rwneg62_2 in62 sn2 3183.098862
Rwneg62_3 in62 sn3 11140.846016
Rwneg62_4 in62 sn4 3183.098862
Rwneg62_5 in62 sn5 11140.846016
Rwneg62_6 in62 sn6 3183.098862
Rwneg62_7 in62 sn7 3183.098862
Rwneg62_8 in62 sn8 11140.846016
Rwneg62_9 in62 sn9 11140.846016
Rwneg62_10 in62 sn10 11140.846016
Rwneg62_11 in62 sn11 11140.846016
Rwneg62_12 in62 sn12 11140.846016
Rwneg62_13 in62 sn13 11140.846016
Rwneg62_14 in62 sn14 11140.846016
Rwneg62_15 in62 sn15 3183.098862
Rwneg62_16 in62 sn16 11140.846016
Rwneg62_17 in62 sn17 3183.098862
Rwneg62_18 in62 sn18 11140.846016
Rwneg62_19 in62 sn19 11140.846016
Rwneg62_20 in62 sn20 3183.098862
Rwneg62_21 in62 sn21 11140.846016
Rwneg62_22 in62 sn22 3183.098862
Rwneg62_23 in62 sn23 11140.846016
Rwneg62_24 in62 sn24 11140.846016
Rwneg62_25 in62 sn25 3183.098862
Rwneg62_26 in62 sn26 3183.098862
Rwneg62_27 in62 sn27 11140.846016
Rwneg62_28 in62 sn28 3183.098862
Rwneg62_29 in62 sn29 11140.846016
Rwneg62_30 in62 sn30 11140.846016
Rwneg62_31 in62 sn31 3183.098862
Rwneg62_32 in62 sn32 3183.098862
Rwneg62_33 in62 sn33 3183.098862
Rwneg62_34 in62 sn34 3183.098862
Rwneg62_35 in62 sn35 11140.846016
Rwneg62_36 in62 sn36 3183.098862
Rwneg62_37 in62 sn37 11140.846016
Rwneg62_38 in62 sn38 11140.846016
Rwneg62_39 in62 sn39 3183.098862
Rwneg62_40 in62 sn40 11140.846016
Rwneg62_41 in62 sn41 11140.846016
Rwneg62_42 in62 sn42 11140.846016
Rwneg62_43 in62 sn43 11140.846016
Rwneg62_44 in62 sn44 11140.846016
Rwneg62_45 in62 sn45 11140.846016
Rwneg62_46 in62 sn46 3183.098862
Rwneg62_47 in62 sn47 3183.098862
Rwneg62_48 in62 sn48 11140.846016
Rwneg62_49 in62 sn49 11140.846016
Rwneg62_50 in62 sn50 11140.846016
Rwneg62_51 in62 sn51 11140.846016
Rwneg62_52 in62 sn52 3183.098862
Rwneg62_53 in62 sn53 11140.846016
Rwneg62_54 in62 sn54 11140.846016
Rwneg62_55 in62 sn55 11140.846016
Rwneg62_56 in62 sn56 3183.098862
Rwneg62_57 in62 sn57 11140.846016
Rwneg62_58 in62 sn58 11140.846016
Rwneg62_59 in62 sn59 11140.846016
Rwneg62_60 in62 sn60 3183.098862
Rwneg62_61 in62 sn61 11140.846016
Rwneg62_62 in62 sn62 3183.098862
Rwneg62_63 in62 sn63 3183.098862
Rwneg62_64 in62 sn64 11140.846016
Rwneg62_65 in62 sn65 11140.846016
Rwneg62_66 in62 sn66 3183.098862
Rwneg62_67 in62 sn67 11140.846016
Rwneg62_68 in62 sn68 11140.846016
Rwneg62_69 in62 sn69 3183.098862
Rwneg62_70 in62 sn70 3183.098862
Rwneg62_71 in62 sn71 11140.846016
Rwneg62_72 in62 sn72 3183.098862
Rwneg62_73 in62 sn73 11140.846016
Rwneg62_74 in62 sn74 11140.846016
Rwneg62_75 in62 sn75 3183.098862
Rwneg62_76 in62 sn76 11140.846016
Rwneg62_77 in62 sn77 11140.846016
Rwneg62_78 in62 sn78 3183.098862
Rwneg62_79 in62 sn79 11140.846016
Rwneg62_80 in62 sn80 3183.098862
Rwneg62_81 in62 sn81 3183.098862
Rwneg62_82 in62 sn82 3183.098862
Rwneg62_83 in62 sn83 11140.846016
Rwneg62_84 in62 sn84 11140.846016
Rwneg62_85 in62 sn85 3183.098862
Rwneg62_86 in62 sn86 3183.098862
Rwneg62_87 in62 sn87 11140.846016
Rwneg62_88 in62 sn88 11140.846016
Rwneg62_89 in62 sn89 11140.846016
Rwneg62_90 in62 sn90 11140.846016
Rwneg62_91 in62 sn91 3183.098862
Rwneg62_92 in62 sn92 3183.098862
Rwneg62_93 in62 sn93 11140.846016
Rwneg62_94 in62 sn94 11140.846016
Rwneg62_95 in62 sn95 3183.098862
Rwneg62_96 in62 sn96 11140.846016
Rwneg62_97 in62 sn97 3183.098862
Rwneg62_98 in62 sn98 3183.098862
Rwneg62_99 in62 sn99 11140.846016
Rwneg62_100 in62 sn100 11140.846016
Rwneg63_1 in63 sn1 11140.846016
Rwneg63_2 in63 sn2 3183.098862
Rwneg63_3 in63 sn3 11140.846016
Rwneg63_4 in63 sn4 3183.098862
Rwneg63_5 in63 sn5 11140.846016
Rwneg63_6 in63 sn6 11140.846016
Rwneg63_7 in63 sn7 3183.098862
Rwneg63_8 in63 sn8 3183.098862
Rwneg63_9 in63 sn9 3183.098862
Rwneg63_10 in63 sn10 11140.846016
Rwneg63_11 in63 sn11 3183.098862
Rwneg63_12 in63 sn12 11140.846016
Rwneg63_13 in63 sn13 11140.846016
Rwneg63_14 in63 sn14 11140.846016
Rwneg63_15 in63 sn15 11140.846016
Rwneg63_16 in63 sn16 11140.846016
Rwneg63_17 in63 sn17 3183.098862
Rwneg63_18 in63 sn18 3183.098862
Rwneg63_19 in63 sn19 11140.846016
Rwneg63_20 in63 sn20 3183.098862
Rwneg63_21 in63 sn21 11140.846016
Rwneg63_22 in63 sn22 11140.846016
Rwneg63_23 in63 sn23 11140.846016
Rwneg63_24 in63 sn24 3183.098862
Rwneg63_25 in63 sn25 11140.846016
Rwneg63_26 in63 sn26 3183.098862
Rwneg63_27 in63 sn27 3183.098862
Rwneg63_28 in63 sn28 11140.846016
Rwneg63_29 in63 sn29 11140.846016
Rwneg63_30 in63 sn30 11140.846016
Rwneg63_31 in63 sn31 3183.098862
Rwneg63_32 in63 sn32 3183.098862
Rwneg63_33 in63 sn33 3183.098862
Rwneg63_34 in63 sn34 11140.846016
Rwneg63_35 in63 sn35 11140.846016
Rwneg63_36 in63 sn36 11140.846016
Rwneg63_37 in63 sn37 3183.098862
Rwneg63_38 in63 sn38 11140.846016
Rwneg63_39 in63 sn39 3183.098862
Rwneg63_40 in63 sn40 11140.846016
Rwneg63_41 in63 sn41 3183.098862
Rwneg63_42 in63 sn42 3183.098862
Rwneg63_43 in63 sn43 3183.098862
Rwneg63_44 in63 sn44 11140.846016
Rwneg63_45 in63 sn45 3183.098862
Rwneg63_46 in63 sn46 3183.098862
Rwneg63_47 in63 sn47 3183.098862
Rwneg63_48 in63 sn48 11140.846016
Rwneg63_49 in63 sn49 11140.846016
Rwneg63_50 in63 sn50 11140.846016
Rwneg63_51 in63 sn51 11140.846016
Rwneg63_52 in63 sn52 3183.098862
Rwneg63_53 in63 sn53 11140.846016
Rwneg63_54 in63 sn54 11140.846016
Rwneg63_55 in63 sn55 3183.098862
Rwneg63_56 in63 sn56 3183.098862
Rwneg63_57 in63 sn57 11140.846016
Rwneg63_58 in63 sn58 11140.846016
Rwneg63_59 in63 sn59 11140.846016
Rwneg63_60 in63 sn60 3183.098862
Rwneg63_61 in63 sn61 3183.098862
Rwneg63_62 in63 sn62 11140.846016
Rwneg63_63 in63 sn63 3183.098862
Rwneg63_64 in63 sn64 3183.098862
Rwneg63_65 in63 sn65 3183.098862
Rwneg63_66 in63 sn66 3183.098862
Rwneg63_67 in63 sn67 3183.098862
Rwneg63_68 in63 sn68 11140.846016
Rwneg63_69 in63 sn69 3183.098862
Rwneg63_70 in63 sn70 3183.098862
Rwneg63_71 in63 sn71 11140.846016
Rwneg63_72 in63 sn72 11140.846016
Rwneg63_73 in63 sn73 11140.846016
Rwneg63_74 in63 sn74 11140.846016
Rwneg63_75 in63 sn75 11140.846016
Rwneg63_76 in63 sn76 11140.846016
Rwneg63_77 in63 sn77 11140.846016
Rwneg63_78 in63 sn78 3183.098862
Rwneg63_79 in63 sn79 11140.846016
Rwneg63_80 in63 sn80 11140.846016
Rwneg63_81 in63 sn81 3183.098862
Rwneg63_82 in63 sn82 11140.846016
Rwneg63_83 in63 sn83 11140.846016
Rwneg63_84 in63 sn84 11140.846016
Rwneg63_85 in63 sn85 11140.846016
Rwneg63_86 in63 sn86 3183.098862
Rwneg63_87 in63 sn87 11140.846016
Rwneg63_88 in63 sn88 11140.846016
Rwneg63_89 in63 sn89 11140.846016
Rwneg63_90 in63 sn90 3183.098862
Rwneg63_91 in63 sn91 3183.098862
Rwneg63_92 in63 sn92 11140.846016
Rwneg63_93 in63 sn93 11140.846016
Rwneg63_94 in63 sn94 11140.846016
Rwneg63_95 in63 sn95 3183.098862
Rwneg63_96 in63 sn96 3183.098862
Rwneg63_97 in63 sn97 11140.846016
Rwneg63_98 in63 sn98 3183.098862
Rwneg63_99 in63 sn99 11140.846016
Rwneg63_100 in63 sn100 11140.846016
Rwneg64_1 in64 sn1 11140.846016
Rwneg64_2 in64 sn2 11140.846016
Rwneg64_3 in64 sn3 11140.846016
Rwneg64_4 in64 sn4 11140.846016
Rwneg64_5 in64 sn5 3183.098862
Rwneg64_6 in64 sn6 11140.846016
Rwneg64_7 in64 sn7 11140.846016
Rwneg64_8 in64 sn8 11140.846016
Rwneg64_9 in64 sn9 3183.098862
Rwneg64_10 in64 sn10 3183.098862
Rwneg64_11 in64 sn11 11140.846016
Rwneg64_12 in64 sn12 3183.098862
Rwneg64_13 in64 sn13 3183.098862
Rwneg64_14 in64 sn14 11140.846016
Rwneg64_15 in64 sn15 3183.098862
Rwneg64_16 in64 sn16 11140.846016
Rwneg64_17 in64 sn17 11140.846016
Rwneg64_18 in64 sn18 3183.098862
Rwneg64_19 in64 sn19 11140.846016
Rwneg64_20 in64 sn20 11140.846016
Rwneg64_21 in64 sn21 11140.846016
Rwneg64_22 in64 sn22 11140.846016
Rwneg64_23 in64 sn23 11140.846016
Rwneg64_24 in64 sn24 11140.846016
Rwneg64_25 in64 sn25 3183.098862
Rwneg64_26 in64 sn26 3183.098862
Rwneg64_27 in64 sn27 3183.098862
Rwneg64_28 in64 sn28 11140.846016
Rwneg64_29 in64 sn29 11140.846016
Rwneg64_30 in64 sn30 3183.098862
Rwneg64_31 in64 sn31 3183.098862
Rwneg64_32 in64 sn32 3183.098862
Rwneg64_33 in64 sn33 3183.098862
Rwneg64_34 in64 sn34 3183.098862
Rwneg64_35 in64 sn35 3183.098862
Rwneg64_36 in64 sn36 3183.098862
Rwneg64_37 in64 sn37 11140.846016
Rwneg64_38 in64 sn38 11140.846016
Rwneg64_39 in64 sn39 11140.846016
Rwneg64_40 in64 sn40 3183.098862
Rwneg64_41 in64 sn41 3183.098862
Rwneg64_42 in64 sn42 11140.846016
Rwneg64_43 in64 sn43 11140.846016
Rwneg64_44 in64 sn44 3183.098862
Rwneg64_45 in64 sn45 11140.846016
Rwneg64_46 in64 sn46 11140.846016
Rwneg64_47 in64 sn47 11140.846016
Rwneg64_48 in64 sn48 3183.098862
Rwneg64_49 in64 sn49 3183.098862
Rwneg64_50 in64 sn50 11140.846016
Rwneg64_51 in64 sn51 11140.846016
Rwneg64_52 in64 sn52 11140.846016
Rwneg64_53 in64 sn53 11140.846016
Rwneg64_54 in64 sn54 3183.098862
Rwneg64_55 in64 sn55 3183.098862
Rwneg64_56 in64 sn56 3183.098862
Rwneg64_57 in64 sn57 3183.098862
Rwneg64_58 in64 sn58 11140.846016
Rwneg64_59 in64 sn59 3183.098862
Rwneg64_60 in64 sn60 3183.098862
Rwneg64_61 in64 sn61 11140.846016
Rwneg64_62 in64 sn62 3183.098862
Rwneg64_63 in64 sn63 3183.098862
Rwneg64_64 in64 sn64 11140.846016
Rwneg64_65 in64 sn65 11140.846016
Rwneg64_66 in64 sn66 11140.846016
Rwneg64_67 in64 sn67 11140.846016
Rwneg64_68 in64 sn68 11140.846016
Rwneg64_69 in64 sn69 11140.846016
Rwneg64_70 in64 sn70 3183.098862
Rwneg64_71 in64 sn71 11140.846016
Rwneg64_72 in64 sn72 11140.846016
Rwneg64_73 in64 sn73 3183.098862
Rwneg64_74 in64 sn74 11140.846016
Rwneg64_75 in64 sn75 11140.846016
Rwneg64_76 in64 sn76 3183.098862
Rwneg64_77 in64 sn77 3183.098862
Rwneg64_78 in64 sn78 3183.098862
Rwneg64_79 in64 sn79 11140.846016
Rwneg64_80 in64 sn80 3183.098862
Rwneg64_81 in64 sn81 11140.846016
Rwneg64_82 in64 sn82 11140.846016
Rwneg64_83 in64 sn83 11140.846016
Rwneg64_84 in64 sn84 11140.846016
Rwneg64_85 in64 sn85 11140.846016
Rwneg64_86 in64 sn86 3183.098862
Rwneg64_87 in64 sn87 3183.098862
Rwneg64_88 in64 sn88 11140.846016
Rwneg64_89 in64 sn89 11140.846016
Rwneg64_90 in64 sn90 3183.098862
Rwneg64_91 in64 sn91 3183.098862
Rwneg64_92 in64 sn92 3183.098862
Rwneg64_93 in64 sn93 3183.098862
Rwneg64_94 in64 sn94 3183.098862
Rwneg64_95 in64 sn95 11140.846016
Rwneg64_96 in64 sn96 11140.846016
Rwneg64_97 in64 sn97 11140.846016
Rwneg64_98 in64 sn98 11140.846016
Rwneg64_99 in64 sn99 3183.098862
Rwneg64_100 in64 sn100 11140.846016
Rwneg65_1 in65 sn1 11140.846016
Rwneg65_2 in65 sn2 3183.098862
Rwneg65_3 in65 sn3 11140.846016
Rwneg65_4 in65 sn4 11140.846016
Rwneg65_5 in65 sn5 11140.846016
Rwneg65_6 in65 sn6 11140.846016
Rwneg65_7 in65 sn7 3183.098862
Rwneg65_8 in65 sn8 11140.846016
Rwneg65_9 in65 sn9 3183.098862
Rwneg65_10 in65 sn10 3183.098862
Rwneg65_11 in65 sn11 11140.846016
Rwneg65_12 in65 sn12 11140.846016
Rwneg65_13 in65 sn13 11140.846016
Rwneg65_14 in65 sn14 11140.846016
Rwneg65_15 in65 sn15 3183.098862
Rwneg65_16 in65 sn16 11140.846016
Rwneg65_17 in65 sn17 11140.846016
Rwneg65_18 in65 sn18 11140.846016
Rwneg65_19 in65 sn19 11140.846016
Rwneg65_20 in65 sn20 11140.846016
Rwneg65_21 in65 sn21 11140.846016
Rwneg65_22 in65 sn22 3183.098862
Rwneg65_23 in65 sn23 3183.098862
Rwneg65_24 in65 sn24 3183.098862
Rwneg65_25 in65 sn25 3183.098862
Rwneg65_26 in65 sn26 3183.098862
Rwneg65_27 in65 sn27 11140.846016
Rwneg65_28 in65 sn28 11140.846016
Rwneg65_29 in65 sn29 11140.846016
Rwneg65_30 in65 sn30 11140.846016
Rwneg65_31 in65 sn31 11140.846016
Rwneg65_32 in65 sn32 3183.098862
Rwneg65_33 in65 sn33 11140.846016
Rwneg65_34 in65 sn34 11140.846016
Rwneg65_35 in65 sn35 3183.098862
Rwneg65_36 in65 sn36 11140.846016
Rwneg65_37 in65 sn37 11140.846016
Rwneg65_38 in65 sn38 11140.846016
Rwneg65_39 in65 sn39 11140.846016
Rwneg65_40 in65 sn40 11140.846016
Rwneg65_41 in65 sn41 3183.098862
Rwneg65_42 in65 sn42 3183.098862
Rwneg65_43 in65 sn43 11140.846016
Rwneg65_44 in65 sn44 3183.098862
Rwneg65_45 in65 sn45 11140.846016
Rwneg65_46 in65 sn46 11140.846016
Rwneg65_47 in65 sn47 11140.846016
Rwneg65_48 in65 sn48 3183.098862
Rwneg65_49 in65 sn49 11140.846016
Rwneg65_50 in65 sn50 3183.098862
Rwneg65_51 in65 sn51 3183.098862
Rwneg65_52 in65 sn52 11140.846016
Rwneg65_53 in65 sn53 11140.846016
Rwneg65_54 in65 sn54 3183.098862
Rwneg65_55 in65 sn55 11140.846016
Rwneg65_56 in65 sn56 3183.098862
Rwneg65_57 in65 sn57 3183.098862
Rwneg65_58 in65 sn58 3183.098862
Rwneg65_59 in65 sn59 3183.098862
Rwneg65_60 in65 sn60 11140.846016
Rwneg65_61 in65 sn61 3183.098862
Rwneg65_62 in65 sn62 11140.846016
Rwneg65_63 in65 sn63 11140.846016
Rwneg65_64 in65 sn64 3183.098862
Rwneg65_65 in65 sn65 11140.846016
Rwneg65_66 in65 sn66 3183.098862
Rwneg65_67 in65 sn67 11140.846016
Rwneg65_68 in65 sn68 11140.846016
Rwneg65_69 in65 sn69 11140.846016
Rwneg65_70 in65 sn70 3183.098862
Rwneg65_71 in65 sn71 11140.846016
Rwneg65_72 in65 sn72 11140.846016
Rwneg65_73 in65 sn73 11140.846016
Rwneg65_74 in65 sn74 3183.098862
Rwneg65_75 in65 sn75 3183.098862
Rwneg65_76 in65 sn76 11140.846016
Rwneg65_77 in65 sn77 3183.098862
Rwneg65_78 in65 sn78 3183.098862
Rwneg65_79 in65 sn79 11140.846016
Rwneg65_80 in65 sn80 3183.098862
Rwneg65_81 in65 sn81 11140.846016
Rwneg65_82 in65 sn82 3183.098862
Rwneg65_83 in65 sn83 3183.098862
Rwneg65_84 in65 sn84 11140.846016
Rwneg65_85 in65 sn85 11140.846016
Rwneg65_86 in65 sn86 11140.846016
Rwneg65_87 in65 sn87 3183.098862
Rwneg65_88 in65 sn88 11140.846016
Rwneg65_89 in65 sn89 11140.846016
Rwneg65_90 in65 sn90 3183.098862
Rwneg65_91 in65 sn91 3183.098862
Rwneg65_92 in65 sn92 11140.846016
Rwneg65_93 in65 sn93 11140.846016
Rwneg65_94 in65 sn94 3183.098862
Rwneg65_95 in65 sn95 11140.846016
Rwneg65_96 in65 sn96 11140.846016
Rwneg65_97 in65 sn97 11140.846016
Rwneg65_98 in65 sn98 11140.846016
Rwneg65_99 in65 sn99 3183.098862
Rwneg65_100 in65 sn100 11140.846016
Rwneg66_1 in66 sn1 11140.846016
Rwneg66_2 in66 sn2 11140.846016
Rwneg66_3 in66 sn3 3183.098862
Rwneg66_4 in66 sn4 11140.846016
Rwneg66_5 in66 sn5 11140.846016
Rwneg66_6 in66 sn6 11140.846016
Rwneg66_7 in66 sn7 11140.846016
Rwneg66_8 in66 sn8 11140.846016
Rwneg66_9 in66 sn9 11140.846016
Rwneg66_10 in66 sn10 3183.098862
Rwneg66_11 in66 sn11 11140.846016
Rwneg66_12 in66 sn12 11140.846016
Rwneg66_13 in66 sn13 11140.846016
Rwneg66_14 in66 sn14 11140.846016
Rwneg66_15 in66 sn15 3183.098862
Rwneg66_16 in66 sn16 3183.098862
Rwneg66_17 in66 sn17 11140.846016
Rwneg66_18 in66 sn18 3183.098862
Rwneg66_19 in66 sn19 3183.098862
Rwneg66_20 in66 sn20 3183.098862
Rwneg66_21 in66 sn21 11140.846016
Rwneg66_22 in66 sn22 11140.846016
Rwneg66_23 in66 sn23 11140.846016
Rwneg66_24 in66 sn24 11140.846016
Rwneg66_25 in66 sn25 11140.846016
Rwneg66_26 in66 sn26 3183.098862
Rwneg66_27 in66 sn27 11140.846016
Rwneg66_28 in66 sn28 11140.846016
Rwneg66_29 in66 sn29 3183.098862
Rwneg66_30 in66 sn30 3183.098862
Rwneg66_31 in66 sn31 3183.098862
Rwneg66_32 in66 sn32 11140.846016
Rwneg66_33 in66 sn33 11140.846016
Rwneg66_34 in66 sn34 11140.846016
Rwneg66_35 in66 sn35 11140.846016
Rwneg66_36 in66 sn36 3183.098862
Rwneg66_37 in66 sn37 11140.846016
Rwneg66_38 in66 sn38 3183.098862
Rwneg66_39 in66 sn39 11140.846016
Rwneg66_40 in66 sn40 11140.846016
Rwneg66_41 in66 sn41 3183.098862
Rwneg66_42 in66 sn42 11140.846016
Rwneg66_43 in66 sn43 11140.846016
Rwneg66_44 in66 sn44 3183.098862
Rwneg66_45 in66 sn45 3183.098862
Rwneg66_46 in66 sn46 3183.098862
Rwneg66_47 in66 sn47 11140.846016
Rwneg66_48 in66 sn48 11140.846016
Rwneg66_49 in66 sn49 11140.846016
Rwneg66_50 in66 sn50 3183.098862
Rwneg66_51 in66 sn51 11140.846016
Rwneg66_52 in66 sn52 3183.098862
Rwneg66_53 in66 sn53 11140.846016
Rwneg66_54 in66 sn54 11140.846016
Rwneg66_55 in66 sn55 3183.098862
Rwneg66_56 in66 sn56 11140.846016
Rwneg66_57 in66 sn57 11140.846016
Rwneg66_58 in66 sn58 11140.846016
Rwneg66_59 in66 sn59 11140.846016
Rwneg66_60 in66 sn60 11140.846016
Rwneg66_61 in66 sn61 3183.098862
Rwneg66_62 in66 sn62 11140.846016
Rwneg66_63 in66 sn63 3183.098862
Rwneg66_64 in66 sn64 3183.098862
Rwneg66_65 in66 sn65 3183.098862
Rwneg66_66 in66 sn66 3183.098862
Rwneg66_67 in66 sn67 11140.846016
Rwneg66_68 in66 sn68 3183.098862
Rwneg66_69 in66 sn69 11140.846016
Rwneg66_70 in66 sn70 11140.846016
Rwneg66_71 in66 sn71 3183.098862
Rwneg66_72 in66 sn72 11140.846016
Rwneg66_73 in66 sn73 11140.846016
Rwneg66_74 in66 sn74 11140.846016
Rwneg66_75 in66 sn75 11140.846016
Rwneg66_76 in66 sn76 11140.846016
Rwneg66_77 in66 sn77 3183.098862
Rwneg66_78 in66 sn78 3183.098862
Rwneg66_79 in66 sn79 11140.846016
Rwneg66_80 in66 sn80 3183.098862
Rwneg66_81 in66 sn81 11140.846016
Rwneg66_82 in66 sn82 3183.098862
Rwneg66_83 in66 sn83 11140.846016
Rwneg66_84 in66 sn84 3183.098862
Rwneg66_85 in66 sn85 11140.846016
Rwneg66_86 in66 sn86 3183.098862
Rwneg66_87 in66 sn87 3183.098862
Rwneg66_88 in66 sn88 11140.846016
Rwneg66_89 in66 sn89 3183.098862
Rwneg66_90 in66 sn90 11140.846016
Rwneg66_91 in66 sn91 11140.846016
Rwneg66_92 in66 sn92 3183.098862
Rwneg66_93 in66 sn93 3183.098862
Rwneg66_94 in66 sn94 3183.098862
Rwneg66_95 in66 sn95 11140.846016
Rwneg66_96 in66 sn96 3183.098862
Rwneg66_97 in66 sn97 11140.846016
Rwneg66_98 in66 sn98 3183.098862
Rwneg66_99 in66 sn99 11140.846016
Rwneg66_100 in66 sn100 3183.098862
Rwneg67_1 in67 sn1 3183.098862
Rwneg67_2 in67 sn2 3183.098862
Rwneg67_3 in67 sn3 3183.098862
Rwneg67_4 in67 sn4 11140.846016
Rwneg67_5 in67 sn5 11140.846016
Rwneg67_6 in67 sn6 11140.846016
Rwneg67_7 in67 sn7 3183.098862
Rwneg67_8 in67 sn8 11140.846016
Rwneg67_9 in67 sn9 3183.098862
Rwneg67_10 in67 sn10 11140.846016
Rwneg67_11 in67 sn11 3183.098862
Rwneg67_12 in67 sn12 11140.846016
Rwneg67_13 in67 sn13 11140.846016
Rwneg67_14 in67 sn14 3183.098862
Rwneg67_15 in67 sn15 11140.846016
Rwneg67_16 in67 sn16 11140.846016
Rwneg67_17 in67 sn17 11140.846016
Rwneg67_18 in67 sn18 3183.098862
Rwneg67_19 in67 sn19 11140.846016
Rwneg67_20 in67 sn20 3183.098862
Rwneg67_21 in67 sn21 11140.846016
Rwneg67_22 in67 sn22 11140.846016
Rwneg67_23 in67 sn23 3183.098862
Rwneg67_24 in67 sn24 11140.846016
Rwneg67_25 in67 sn25 11140.846016
Rwneg67_26 in67 sn26 11140.846016
Rwneg67_27 in67 sn27 11140.846016
Rwneg67_28 in67 sn28 3183.098862
Rwneg67_29 in67 sn29 11140.846016
Rwneg67_30 in67 sn30 3183.098862
Rwneg67_31 in67 sn31 11140.846016
Rwneg67_32 in67 sn32 11140.846016
Rwneg67_33 in67 sn33 11140.846016
Rwneg67_34 in67 sn34 3183.098862
Rwneg67_35 in67 sn35 11140.846016
Rwneg67_36 in67 sn36 11140.846016
Rwneg67_37 in67 sn37 11140.846016
Rwneg67_38 in67 sn38 11140.846016
Rwneg67_39 in67 sn39 3183.098862
Rwneg67_40 in67 sn40 11140.846016
Rwneg67_41 in67 sn41 11140.846016
Rwneg67_42 in67 sn42 11140.846016
Rwneg67_43 in67 sn43 11140.846016
Rwneg67_44 in67 sn44 11140.846016
Rwneg67_45 in67 sn45 3183.098862
Rwneg67_46 in67 sn46 3183.098862
Rwneg67_47 in67 sn47 3183.098862
Rwneg67_48 in67 sn48 11140.846016
Rwneg67_49 in67 sn49 11140.846016
Rwneg67_50 in67 sn50 3183.098862
Rwneg67_51 in67 sn51 11140.846016
Rwneg67_52 in67 sn52 11140.846016
Rwneg67_53 in67 sn53 11140.846016
Rwneg67_54 in67 sn54 11140.846016
Rwneg67_55 in67 sn55 3183.098862
Rwneg67_56 in67 sn56 3183.098862
Rwneg67_57 in67 sn57 3183.098862
Rwneg67_58 in67 sn58 11140.846016
Rwneg67_59 in67 sn59 3183.098862
Rwneg67_60 in67 sn60 3183.098862
Rwneg67_61 in67 sn61 3183.098862
Rwneg67_62 in67 sn62 3183.098862
Rwneg67_63 in67 sn63 3183.098862
Rwneg67_64 in67 sn64 11140.846016
Rwneg67_65 in67 sn65 3183.098862
Rwneg67_66 in67 sn66 11140.846016
Rwneg67_67 in67 sn67 11140.846016
Rwneg67_68 in67 sn68 11140.846016
Rwneg67_69 in67 sn69 3183.098862
Rwneg67_70 in67 sn70 11140.846016
Rwneg67_71 in67 sn71 3183.098862
Rwneg67_72 in67 sn72 11140.846016
Rwneg67_73 in67 sn73 3183.098862
Rwneg67_74 in67 sn74 11140.846016
Rwneg67_75 in67 sn75 11140.846016
Rwneg67_76 in67 sn76 11140.846016
Rwneg67_77 in67 sn77 3183.098862
Rwneg67_78 in67 sn78 11140.846016
Rwneg67_79 in67 sn79 3183.098862
Rwneg67_80 in67 sn80 11140.846016
Rwneg67_81 in67 sn81 11140.846016
Rwneg67_82 in67 sn82 3183.098862
Rwneg67_83 in67 sn83 3183.098862
Rwneg67_84 in67 sn84 11140.846016
Rwneg67_85 in67 sn85 11140.846016
Rwneg67_86 in67 sn86 3183.098862
Rwneg67_87 in67 sn87 11140.846016
Rwneg67_88 in67 sn88 3183.098862
Rwneg67_89 in67 sn89 3183.098862
Rwneg67_90 in67 sn90 3183.098862
Rwneg67_91 in67 sn91 11140.846016
Rwneg67_92 in67 sn92 11140.846016
Rwneg67_93 in67 sn93 3183.098862
Rwneg67_94 in67 sn94 11140.846016
Rwneg67_95 in67 sn95 3183.098862
Rwneg67_96 in67 sn96 11140.846016
Rwneg67_97 in67 sn97 11140.846016
Rwneg67_98 in67 sn98 3183.098862
Rwneg67_99 in67 sn99 11140.846016
Rwneg67_100 in67 sn100 11140.846016
Rwneg68_1 in68 sn1 3183.098862
Rwneg68_2 in68 sn2 11140.846016
Rwneg68_3 in68 sn3 11140.846016
Rwneg68_4 in68 sn4 11140.846016
Rwneg68_5 in68 sn5 11140.846016
Rwneg68_6 in68 sn6 3183.098862
Rwneg68_7 in68 sn7 3183.098862
Rwneg68_8 in68 sn8 11140.846016
Rwneg68_9 in68 sn9 3183.098862
Rwneg68_10 in68 sn10 11140.846016
Rwneg68_11 in68 sn11 3183.098862
Rwneg68_12 in68 sn12 3183.098862
Rwneg68_13 in68 sn13 11140.846016
Rwneg68_14 in68 sn14 3183.098862
Rwneg68_15 in68 sn15 11140.846016
Rwneg68_16 in68 sn16 11140.846016
Rwneg68_17 in68 sn17 11140.846016
Rwneg68_18 in68 sn18 11140.846016
Rwneg68_19 in68 sn19 3183.098862
Rwneg68_20 in68 sn20 3183.098862
Rwneg68_21 in68 sn21 3183.098862
Rwneg68_22 in68 sn22 11140.846016
Rwneg68_23 in68 sn23 11140.846016
Rwneg68_24 in68 sn24 3183.098862
Rwneg68_25 in68 sn25 11140.846016
Rwneg68_26 in68 sn26 3183.098862
Rwneg68_27 in68 sn27 3183.098862
Rwneg68_28 in68 sn28 3183.098862
Rwneg68_29 in68 sn29 11140.846016
Rwneg68_30 in68 sn30 11140.846016
Rwneg68_31 in68 sn31 3183.098862
Rwneg68_32 in68 sn32 11140.846016
Rwneg68_33 in68 sn33 11140.846016
Rwneg68_34 in68 sn34 3183.098862
Rwneg68_35 in68 sn35 3183.098862
Rwneg68_36 in68 sn36 11140.846016
Rwneg68_37 in68 sn37 11140.846016
Rwneg68_38 in68 sn38 3183.098862
Rwneg68_39 in68 sn39 11140.846016
Rwneg68_40 in68 sn40 11140.846016
Rwneg68_41 in68 sn41 3183.098862
Rwneg68_42 in68 sn42 11140.846016
Rwneg68_43 in68 sn43 3183.098862
Rwneg68_44 in68 sn44 11140.846016
Rwneg68_45 in68 sn45 11140.846016
Rwneg68_46 in68 sn46 11140.846016
Rwneg68_47 in68 sn47 3183.098862
Rwneg68_48 in68 sn48 11140.846016
Rwneg68_49 in68 sn49 11140.846016
Rwneg68_50 in68 sn50 11140.846016
Rwneg68_51 in68 sn51 3183.098862
Rwneg68_52 in68 sn52 3183.098862
Rwneg68_53 in68 sn53 11140.846016
Rwneg68_54 in68 sn54 11140.846016
Rwneg68_55 in68 sn55 3183.098862
Rwneg68_56 in68 sn56 11140.846016
Rwneg68_57 in68 sn57 11140.846016
Rwneg68_58 in68 sn58 11140.846016
Rwneg68_59 in68 sn59 11140.846016
Rwneg68_60 in68 sn60 3183.098862
Rwneg68_61 in68 sn61 11140.846016
Rwneg68_62 in68 sn62 3183.098862
Rwneg68_63 in68 sn63 3183.098862
Rwneg68_64 in68 sn64 3183.098862
Rwneg68_65 in68 sn65 11140.846016
Rwneg68_66 in68 sn66 3183.098862
Rwneg68_67 in68 sn67 11140.846016
Rwneg68_68 in68 sn68 3183.098862
Rwneg68_69 in68 sn69 3183.098862
Rwneg68_70 in68 sn70 11140.846016
Rwneg68_71 in68 sn71 3183.098862
Rwneg68_72 in68 sn72 11140.846016
Rwneg68_73 in68 sn73 11140.846016
Rwneg68_74 in68 sn74 3183.098862
Rwneg68_75 in68 sn75 3183.098862
Rwneg68_76 in68 sn76 11140.846016
Rwneg68_77 in68 sn77 3183.098862
Rwneg68_78 in68 sn78 3183.098862
Rwneg68_79 in68 sn79 3183.098862
Rwneg68_80 in68 sn80 11140.846016
Rwneg68_81 in68 sn81 11140.846016
Rwneg68_82 in68 sn82 11140.846016
Rwneg68_83 in68 sn83 3183.098862
Rwneg68_84 in68 sn84 11140.846016
Rwneg68_85 in68 sn85 11140.846016
Rwneg68_86 in68 sn86 11140.846016
Rwneg68_87 in68 sn87 11140.846016
Rwneg68_88 in68 sn88 11140.846016
Rwneg68_89 in68 sn89 11140.846016
Rwneg68_90 in68 sn90 3183.098862
Rwneg68_91 in68 sn91 3183.098862
Rwneg68_92 in68 sn92 3183.098862
Rwneg68_93 in68 sn93 3183.098862
Rwneg68_94 in68 sn94 11140.846016
Rwneg68_95 in68 sn95 3183.098862
Rwneg68_96 in68 sn96 11140.846016
Rwneg68_97 in68 sn97 11140.846016
Rwneg68_98 in68 sn98 3183.098862
Rwneg68_99 in68 sn99 3183.098862
Rwneg68_100 in68 sn100 3183.098862
Rwneg69_1 in69 sn1 11140.846016
Rwneg69_2 in69 sn2 11140.846016
Rwneg69_3 in69 sn3 3183.098862
Rwneg69_4 in69 sn4 11140.846016
Rwneg69_5 in69 sn5 11140.846016
Rwneg69_6 in69 sn6 11140.846016
Rwneg69_7 in69 sn7 11140.846016
Rwneg69_8 in69 sn8 11140.846016
Rwneg69_9 in69 sn9 3183.098862
Rwneg69_10 in69 sn10 3183.098862
Rwneg69_11 in69 sn11 11140.846016
Rwneg69_12 in69 sn12 3183.098862
Rwneg69_13 in69 sn13 11140.846016
Rwneg69_14 in69 sn14 11140.846016
Rwneg69_15 in69 sn15 11140.846016
Rwneg69_16 in69 sn16 11140.846016
Rwneg69_17 in69 sn17 11140.846016
Rwneg69_18 in69 sn18 3183.098862
Rwneg69_19 in69 sn19 11140.846016
Rwneg69_20 in69 sn20 11140.846016
Rwneg69_21 in69 sn21 3183.098862
Rwneg69_22 in69 sn22 11140.846016
Rwneg69_23 in69 sn23 11140.846016
Rwneg69_24 in69 sn24 3183.098862
Rwneg69_25 in69 sn25 3183.098862
Rwneg69_26 in69 sn26 3183.098862
Rwneg69_27 in69 sn27 11140.846016
Rwneg69_28 in69 sn28 3183.098862
Rwneg69_29 in69 sn29 11140.846016
Rwneg69_30 in69 sn30 11140.846016
Rwneg69_31 in69 sn31 11140.846016
Rwneg69_32 in69 sn32 11140.846016
Rwneg69_33 in69 sn33 11140.846016
Rwneg69_34 in69 sn34 3183.098862
Rwneg69_35 in69 sn35 3183.098862
Rwneg69_36 in69 sn36 11140.846016
Rwneg69_37 in69 sn37 11140.846016
Rwneg69_38 in69 sn38 11140.846016
Rwneg69_39 in69 sn39 11140.846016
Rwneg69_40 in69 sn40 3183.098862
Rwneg69_41 in69 sn41 3183.098862
Rwneg69_42 in69 sn42 3183.098862
Rwneg69_43 in69 sn43 11140.846016
Rwneg69_44 in69 sn44 3183.098862
Rwneg69_45 in69 sn45 11140.846016
Rwneg69_46 in69 sn46 11140.846016
Rwneg69_47 in69 sn47 11140.846016
Rwneg69_48 in69 sn48 11140.846016
Rwneg69_49 in69 sn49 11140.846016
Rwneg69_50 in69 sn50 3183.098862
Rwneg69_51 in69 sn51 11140.846016
Rwneg69_52 in69 sn52 11140.846016
Rwneg69_53 in69 sn53 11140.846016
Rwneg69_54 in69 sn54 3183.098862
Rwneg69_55 in69 sn55 3183.098862
Rwneg69_56 in69 sn56 3183.098862
Rwneg69_57 in69 sn57 11140.846016
Rwneg69_58 in69 sn58 3183.098862
Rwneg69_59 in69 sn59 3183.098862
Rwneg69_60 in69 sn60 3183.098862
Rwneg69_61 in69 sn61 11140.846016
Rwneg69_62 in69 sn62 11140.846016
Rwneg69_63 in69 sn63 11140.846016
Rwneg69_64 in69 sn64 11140.846016
Rwneg69_65 in69 sn65 11140.846016
Rwneg69_66 in69 sn66 11140.846016
Rwneg69_67 in69 sn67 3183.098862
Rwneg69_68 in69 sn68 11140.846016
Rwneg69_69 in69 sn69 11140.846016
Rwneg69_70 in69 sn70 11140.846016
Rwneg69_71 in69 sn71 11140.846016
Rwneg69_72 in69 sn72 3183.098862
Rwneg69_73 in69 sn73 3183.098862
Rwneg69_74 in69 sn74 3183.098862
Rwneg69_75 in69 sn75 3183.098862
Rwneg69_76 in69 sn76 3183.098862
Rwneg69_77 in69 sn77 3183.098862
Rwneg69_78 in69 sn78 11140.846016
Rwneg69_79 in69 sn79 3183.098862
Rwneg69_80 in69 sn80 3183.098862
Rwneg69_81 in69 sn81 11140.846016
Rwneg69_82 in69 sn82 3183.098862
Rwneg69_83 in69 sn83 3183.098862
Rwneg69_84 in69 sn84 11140.846016
Rwneg69_85 in69 sn85 11140.846016
Rwneg69_86 in69 sn86 3183.098862
Rwneg69_87 in69 sn87 3183.098862
Rwneg69_88 in69 sn88 11140.846016
Rwneg69_89 in69 sn89 3183.098862
Rwneg69_90 in69 sn90 3183.098862
Rwneg69_91 in69 sn91 11140.846016
Rwneg69_92 in69 sn92 3183.098862
Rwneg69_93 in69 sn93 11140.846016
Rwneg69_94 in69 sn94 11140.846016
Rwneg69_95 in69 sn95 11140.846016
Rwneg69_96 in69 sn96 3183.098862
Rwneg69_97 in69 sn97 3183.098862
Rwneg69_98 in69 sn98 3183.098862
Rwneg69_99 in69 sn99 3183.098862
Rwneg69_100 in69 sn100 11140.846016
Rwneg70_1 in70 sn1 11140.846016
Rwneg70_2 in70 sn2 11140.846016
Rwneg70_3 in70 sn3 11140.846016
Rwneg70_4 in70 sn4 3183.098862
Rwneg70_5 in70 sn5 3183.098862
Rwneg70_6 in70 sn6 3183.098862
Rwneg70_7 in70 sn7 3183.098862
Rwneg70_8 in70 sn8 3183.098862
Rwneg70_9 in70 sn9 3183.098862
Rwneg70_10 in70 sn10 11140.846016
Rwneg70_11 in70 sn11 11140.846016
Rwneg70_12 in70 sn12 3183.098862
Rwneg70_13 in70 sn13 11140.846016
Rwneg70_14 in70 sn14 3183.098862
Rwneg70_15 in70 sn15 3183.098862
Rwneg70_16 in70 sn16 11140.846016
Rwneg70_17 in70 sn17 11140.846016
Rwneg70_18 in70 sn18 3183.098862
Rwneg70_19 in70 sn19 3183.098862
Rwneg70_20 in70 sn20 11140.846016
Rwneg70_21 in70 sn21 11140.846016
Rwneg70_22 in70 sn22 3183.098862
Rwneg70_23 in70 sn23 11140.846016
Rwneg70_24 in70 sn24 11140.846016
Rwneg70_25 in70 sn25 3183.098862
Rwneg70_26 in70 sn26 3183.098862
Rwneg70_27 in70 sn27 11140.846016
Rwneg70_28 in70 sn28 3183.098862
Rwneg70_29 in70 sn29 11140.846016
Rwneg70_30 in70 sn30 3183.098862
Rwneg70_31 in70 sn31 3183.098862
Rwneg70_32 in70 sn32 3183.098862
Rwneg70_33 in70 sn33 11140.846016
Rwneg70_34 in70 sn34 11140.846016
Rwneg70_35 in70 sn35 3183.098862
Rwneg70_36 in70 sn36 3183.098862
Rwneg70_37 in70 sn37 11140.846016
Rwneg70_38 in70 sn38 11140.846016
Rwneg70_39 in70 sn39 3183.098862
Rwneg70_40 in70 sn40 11140.846016
Rwneg70_41 in70 sn41 3183.098862
Rwneg70_42 in70 sn42 3183.098862
Rwneg70_43 in70 sn43 11140.846016
Rwneg70_44 in70 sn44 3183.098862
Rwneg70_45 in70 sn45 11140.846016
Rwneg70_46 in70 sn46 3183.098862
Rwneg70_47 in70 sn47 11140.846016
Rwneg70_48 in70 sn48 3183.098862
Rwneg70_49 in70 sn49 11140.846016
Rwneg70_50 in70 sn50 3183.098862
Rwneg70_51 in70 sn51 11140.846016
Rwneg70_52 in70 sn52 11140.846016
Rwneg70_53 in70 sn53 11140.846016
Rwneg70_54 in70 sn54 3183.098862
Rwneg70_55 in70 sn55 3183.098862
Rwneg70_56 in70 sn56 11140.846016
Rwneg70_57 in70 sn57 11140.846016
Rwneg70_58 in70 sn58 3183.098862
Rwneg70_59 in70 sn59 11140.846016
Rwneg70_60 in70 sn60 3183.098862
Rwneg70_61 in70 sn61 3183.098862
Rwneg70_62 in70 sn62 3183.098862
Rwneg70_63 in70 sn63 3183.098862
Rwneg70_64 in70 sn64 11140.846016
Rwneg70_65 in70 sn65 11140.846016
Rwneg70_66 in70 sn66 3183.098862
Rwneg70_67 in70 sn67 3183.098862
Rwneg70_68 in70 sn68 3183.098862
Rwneg70_69 in70 sn69 11140.846016
Rwneg70_70 in70 sn70 3183.098862
Rwneg70_71 in70 sn71 11140.846016
Rwneg70_72 in70 sn72 11140.846016
Rwneg70_73 in70 sn73 11140.846016
Rwneg70_74 in70 sn74 3183.098862
Rwneg70_75 in70 sn75 11140.846016
Rwneg70_76 in70 sn76 11140.846016
Rwneg70_77 in70 sn77 3183.098862
Rwneg70_78 in70 sn78 3183.098862
Rwneg70_79 in70 sn79 3183.098862
Rwneg70_80 in70 sn80 11140.846016
Rwneg70_81 in70 sn81 3183.098862
Rwneg70_82 in70 sn82 3183.098862
Rwneg70_83 in70 sn83 11140.846016
Rwneg70_84 in70 sn84 3183.098862
Rwneg70_85 in70 sn85 11140.846016
Rwneg70_86 in70 sn86 3183.098862
Rwneg70_87 in70 sn87 3183.098862
Rwneg70_88 in70 sn88 11140.846016
Rwneg70_89 in70 sn89 11140.846016
Rwneg70_90 in70 sn90 3183.098862
Rwneg70_91 in70 sn91 11140.846016
Rwneg70_92 in70 sn92 3183.098862
Rwneg70_93 in70 sn93 3183.098862
Rwneg70_94 in70 sn94 11140.846016
Rwneg70_95 in70 sn95 3183.098862
Rwneg70_96 in70 sn96 11140.846016
Rwneg70_97 in70 sn97 11140.846016
Rwneg70_98 in70 sn98 3183.098862
Rwneg70_99 in70 sn99 11140.846016
Rwneg70_100 in70 sn100 3183.098862
Rwneg71_1 in71 sn1 11140.846016
Rwneg71_2 in71 sn2 3183.098862
Rwneg71_3 in71 sn3 11140.846016
Rwneg71_4 in71 sn4 11140.846016
Rwneg71_5 in71 sn5 11140.846016
Rwneg71_6 in71 sn6 11140.846016
Rwneg71_7 in71 sn7 3183.098862
Rwneg71_8 in71 sn8 11140.846016
Rwneg71_9 in71 sn9 3183.098862
Rwneg71_10 in71 sn10 3183.098862
Rwneg71_11 in71 sn11 11140.846016
Rwneg71_12 in71 sn12 3183.098862
Rwneg71_13 in71 sn13 11140.846016
Rwneg71_14 in71 sn14 3183.098862
Rwneg71_15 in71 sn15 3183.098862
Rwneg71_16 in71 sn16 3183.098862
Rwneg71_17 in71 sn17 11140.846016
Rwneg71_18 in71 sn18 11140.846016
Rwneg71_19 in71 sn19 11140.846016
Rwneg71_20 in71 sn20 3183.098862
Rwneg71_21 in71 sn21 11140.846016
Rwneg71_22 in71 sn22 11140.846016
Rwneg71_23 in71 sn23 11140.846016
Rwneg71_24 in71 sn24 11140.846016
Rwneg71_25 in71 sn25 3183.098862
Rwneg71_26 in71 sn26 11140.846016
Rwneg71_27 in71 sn27 3183.098862
Rwneg71_28 in71 sn28 3183.098862
Rwneg71_29 in71 sn29 11140.846016
Rwneg71_30 in71 sn30 3183.098862
Rwneg71_31 in71 sn31 11140.846016
Rwneg71_32 in71 sn32 3183.098862
Rwneg71_33 in71 sn33 11140.846016
Rwneg71_34 in71 sn34 3183.098862
Rwneg71_35 in71 sn35 11140.846016
Rwneg71_36 in71 sn36 3183.098862
Rwneg71_37 in71 sn37 11140.846016
Rwneg71_38 in71 sn38 11140.846016
Rwneg71_39 in71 sn39 3183.098862
Rwneg71_40 in71 sn40 3183.098862
Rwneg71_41 in71 sn41 3183.098862
Rwneg71_42 in71 sn42 3183.098862
Rwneg71_43 in71 sn43 11140.846016
Rwneg71_44 in71 sn44 3183.098862
Rwneg71_45 in71 sn45 11140.846016
Rwneg71_46 in71 sn46 3183.098862
Rwneg71_47 in71 sn47 11140.846016
Rwneg71_48 in71 sn48 3183.098862
Rwneg71_49 in71 sn49 11140.846016
Rwneg71_50 in71 sn50 3183.098862
Rwneg71_51 in71 sn51 11140.846016
Rwneg71_52 in71 sn52 11140.846016
Rwneg71_53 in71 sn53 11140.846016
Rwneg71_54 in71 sn54 11140.846016
Rwneg71_55 in71 sn55 11140.846016
Rwneg71_56 in71 sn56 11140.846016
Rwneg71_57 in71 sn57 3183.098862
Rwneg71_58 in71 sn58 11140.846016
Rwneg71_59 in71 sn59 11140.846016
Rwneg71_60 in71 sn60 11140.846016
Rwneg71_61 in71 sn61 3183.098862
Rwneg71_62 in71 sn62 3183.098862
Rwneg71_63 in71 sn63 3183.098862
Rwneg71_64 in71 sn64 11140.846016
Rwneg71_65 in71 sn65 3183.098862
Rwneg71_66 in71 sn66 3183.098862
Rwneg71_67 in71 sn67 11140.846016
Rwneg71_68 in71 sn68 11140.846016
Rwneg71_69 in71 sn69 11140.846016
Rwneg71_70 in71 sn70 11140.846016
Rwneg71_71 in71 sn71 3183.098862
Rwneg71_72 in71 sn72 3183.098862
Rwneg71_73 in71 sn73 3183.098862
Rwneg71_74 in71 sn74 3183.098862
Rwneg71_75 in71 sn75 11140.846016
Rwneg71_76 in71 sn76 3183.098862
Rwneg71_77 in71 sn77 3183.098862
Rwneg71_78 in71 sn78 3183.098862
Rwneg71_79 in71 sn79 11140.846016
Rwneg71_80 in71 sn80 11140.846016
Rwneg71_81 in71 sn81 3183.098862
Rwneg71_82 in71 sn82 3183.098862
Rwneg71_83 in71 sn83 11140.846016
Rwneg71_84 in71 sn84 3183.098862
Rwneg71_85 in71 sn85 11140.846016
Rwneg71_86 in71 sn86 11140.846016
Rwneg71_87 in71 sn87 3183.098862
Rwneg71_88 in71 sn88 11140.846016
Rwneg71_89 in71 sn89 11140.846016
Rwneg71_90 in71 sn90 3183.098862
Rwneg71_91 in71 sn91 11140.846016
Rwneg71_92 in71 sn92 3183.098862
Rwneg71_93 in71 sn93 3183.098862
Rwneg71_94 in71 sn94 3183.098862
Rwneg71_95 in71 sn95 11140.846016
Rwneg71_96 in71 sn96 11140.846016
Rwneg71_97 in71 sn97 3183.098862
Rwneg71_98 in71 sn98 3183.098862
Rwneg71_99 in71 sn99 11140.846016
Rwneg71_100 in71 sn100 3183.098862
Rwneg72_1 in72 sn1 11140.846016
Rwneg72_2 in72 sn2 11140.846016
Rwneg72_3 in72 sn3 3183.098862
Rwneg72_4 in72 sn4 3183.098862
Rwneg72_5 in72 sn5 11140.846016
Rwneg72_6 in72 sn6 11140.846016
Rwneg72_7 in72 sn7 11140.846016
Rwneg72_8 in72 sn8 11140.846016
Rwneg72_9 in72 sn9 11140.846016
Rwneg72_10 in72 sn10 3183.098862
Rwneg72_11 in72 sn11 3183.098862
Rwneg72_12 in72 sn12 3183.098862
Rwneg72_13 in72 sn13 11140.846016
Rwneg72_14 in72 sn14 3183.098862
Rwneg72_15 in72 sn15 11140.846016
Rwneg72_16 in72 sn16 11140.846016
Rwneg72_17 in72 sn17 11140.846016
Rwneg72_18 in72 sn18 11140.846016
Rwneg72_19 in72 sn19 3183.098862
Rwneg72_20 in72 sn20 3183.098862
Rwneg72_21 in72 sn21 11140.846016
Rwneg72_22 in72 sn22 11140.846016
Rwneg72_23 in72 sn23 11140.846016
Rwneg72_24 in72 sn24 11140.846016
Rwneg72_25 in72 sn25 11140.846016
Rwneg72_26 in72 sn26 3183.098862
Rwneg72_27 in72 sn27 3183.098862
Rwneg72_28 in72 sn28 11140.846016
Rwneg72_29 in72 sn29 3183.098862
Rwneg72_30 in72 sn30 3183.098862
Rwneg72_31 in72 sn31 11140.846016
Rwneg72_32 in72 sn32 3183.098862
Rwneg72_33 in72 sn33 3183.098862
Rwneg72_34 in72 sn34 11140.846016
Rwneg72_35 in72 sn35 11140.846016
Rwneg72_36 in72 sn36 3183.098862
Rwneg72_37 in72 sn37 3183.098862
Rwneg72_38 in72 sn38 3183.098862
Rwneg72_39 in72 sn39 11140.846016
Rwneg72_40 in72 sn40 3183.098862
Rwneg72_41 in72 sn41 3183.098862
Rwneg72_42 in72 sn42 11140.846016
Rwneg72_43 in72 sn43 11140.846016
Rwneg72_44 in72 sn44 11140.846016
Rwneg72_45 in72 sn45 11140.846016
Rwneg72_46 in72 sn46 3183.098862
Rwneg72_47 in72 sn47 3183.098862
Rwneg72_48 in72 sn48 3183.098862
Rwneg72_49 in72 sn49 11140.846016
Rwneg72_50 in72 sn50 11140.846016
Rwneg72_51 in72 sn51 3183.098862
Rwneg72_52 in72 sn52 11140.846016
Rwneg72_53 in72 sn53 3183.098862
Rwneg72_54 in72 sn54 3183.098862
Rwneg72_55 in72 sn55 11140.846016
Rwneg72_56 in72 sn56 11140.846016
Rwneg72_57 in72 sn57 3183.098862
Rwneg72_58 in72 sn58 11140.846016
Rwneg72_59 in72 sn59 11140.846016
Rwneg72_60 in72 sn60 11140.846016
Rwneg72_61 in72 sn61 3183.098862
Rwneg72_62 in72 sn62 3183.098862
Rwneg72_63 in72 sn63 11140.846016
Rwneg72_64 in72 sn64 11140.846016
Rwneg72_65 in72 sn65 3183.098862
Rwneg72_66 in72 sn66 11140.846016
Rwneg72_67 in72 sn67 11140.846016
Rwneg72_68 in72 sn68 11140.846016
Rwneg72_69 in72 sn69 3183.098862
Rwneg72_70 in72 sn70 3183.098862
Rwneg72_71 in72 sn71 3183.098862
Rwneg72_72 in72 sn72 3183.098862
Rwneg72_73 in72 sn73 11140.846016
Rwneg72_74 in72 sn74 3183.098862
Rwneg72_75 in72 sn75 11140.846016
Rwneg72_76 in72 sn76 11140.846016
Rwneg72_77 in72 sn77 3183.098862
Rwneg72_78 in72 sn78 11140.846016
Rwneg72_79 in72 sn79 3183.098862
Rwneg72_80 in72 sn80 3183.098862
Rwneg72_81 in72 sn81 3183.098862
Rwneg72_82 in72 sn82 3183.098862
Rwneg72_83 in72 sn83 3183.098862
Rwneg72_84 in72 sn84 3183.098862
Rwneg72_85 in72 sn85 11140.846016
Rwneg72_86 in72 sn86 3183.098862
Rwneg72_87 in72 sn87 11140.846016
Rwneg72_88 in72 sn88 11140.846016
Rwneg72_89 in72 sn89 11140.846016
Rwneg72_90 in72 sn90 3183.098862
Rwneg72_91 in72 sn91 3183.098862
Rwneg72_92 in72 sn92 3183.098862
Rwneg72_93 in72 sn93 3183.098862
Rwneg72_94 in72 sn94 3183.098862
Rwneg72_95 in72 sn95 11140.846016
Rwneg72_96 in72 sn96 3183.098862
Rwneg72_97 in72 sn97 3183.098862
Rwneg72_98 in72 sn98 11140.846016
Rwneg72_99 in72 sn99 11140.846016
Rwneg72_100 in72 sn100 3183.098862
Rwneg73_1 in73 sn1 3183.098862
Rwneg73_2 in73 sn2 11140.846016
Rwneg73_3 in73 sn3 11140.846016
Rwneg73_4 in73 sn4 3183.098862
Rwneg73_5 in73 sn5 11140.846016
Rwneg73_6 in73 sn6 3183.098862
Rwneg73_7 in73 sn7 3183.098862
Rwneg73_8 in73 sn8 11140.846016
Rwneg73_9 in73 sn9 11140.846016
Rwneg73_10 in73 sn10 11140.846016
Rwneg73_11 in73 sn11 11140.846016
Rwneg73_12 in73 sn12 11140.846016
Rwneg73_13 in73 sn13 11140.846016
Rwneg73_14 in73 sn14 11140.846016
Rwneg73_15 in73 sn15 11140.846016
Rwneg73_16 in73 sn16 11140.846016
Rwneg73_17 in73 sn17 3183.098862
Rwneg73_18 in73 sn18 3183.098862
Rwneg73_19 in73 sn19 11140.846016
Rwneg73_20 in73 sn20 3183.098862
Rwneg73_21 in73 sn21 3183.098862
Rwneg73_22 in73 sn22 11140.846016
Rwneg73_23 in73 sn23 11140.846016
Rwneg73_24 in73 sn24 3183.098862
Rwneg73_25 in73 sn25 3183.098862
Rwneg73_26 in73 sn26 3183.098862
Rwneg73_27 in73 sn27 11140.846016
Rwneg73_28 in73 sn28 11140.846016
Rwneg73_29 in73 sn29 3183.098862
Rwneg73_30 in73 sn30 3183.098862
Rwneg73_31 in73 sn31 11140.846016
Rwneg73_32 in73 sn32 11140.846016
Rwneg73_33 in73 sn33 3183.098862
Rwneg73_34 in73 sn34 3183.098862
Rwneg73_35 in73 sn35 11140.846016
Rwneg73_36 in73 sn36 3183.098862
Rwneg73_37 in73 sn37 11140.846016
Rwneg73_38 in73 sn38 11140.846016
Rwneg73_39 in73 sn39 3183.098862
Rwneg73_40 in73 sn40 3183.098862
Rwneg73_41 in73 sn41 3183.098862
Rwneg73_42 in73 sn42 3183.098862
Rwneg73_43 in73 sn43 3183.098862
Rwneg73_44 in73 sn44 11140.846016
Rwneg73_45 in73 sn45 11140.846016
Rwneg73_46 in73 sn46 3183.098862
Rwneg73_47 in73 sn47 3183.098862
Rwneg73_48 in73 sn48 11140.846016
Rwneg73_49 in73 sn49 3183.098862
Rwneg73_50 in73 sn50 3183.098862
Rwneg73_51 in73 sn51 3183.098862
Rwneg73_52 in73 sn52 11140.846016
Rwneg73_53 in73 sn53 11140.846016
Rwneg73_54 in73 sn54 11140.846016
Rwneg73_55 in73 sn55 11140.846016
Rwneg73_56 in73 sn56 11140.846016
Rwneg73_57 in73 sn57 11140.846016
Rwneg73_58 in73 sn58 11140.846016
Rwneg73_59 in73 sn59 11140.846016
Rwneg73_60 in73 sn60 3183.098862
Rwneg73_61 in73 sn61 11140.846016
Rwneg73_62 in73 sn62 11140.846016
Rwneg73_63 in73 sn63 11140.846016
Rwneg73_64 in73 sn64 11140.846016
Rwneg73_65 in73 sn65 11140.846016
Rwneg73_66 in73 sn66 3183.098862
Rwneg73_67 in73 sn67 11140.846016
Rwneg73_68 in73 sn68 11140.846016
Rwneg73_69 in73 sn69 11140.846016
Rwneg73_70 in73 sn70 11140.846016
Rwneg73_71 in73 sn71 3183.098862
Rwneg73_72 in73 sn72 3183.098862
Rwneg73_73 in73 sn73 11140.846016
Rwneg73_74 in73 sn74 3183.098862
Rwneg73_75 in73 sn75 3183.098862
Rwneg73_76 in73 sn76 3183.098862
Rwneg73_77 in73 sn77 11140.846016
Rwneg73_78 in73 sn78 11140.846016
Rwneg73_79 in73 sn79 3183.098862
Rwneg73_80 in73 sn80 3183.098862
Rwneg73_81 in73 sn81 11140.846016
Rwneg73_82 in73 sn82 11140.846016
Rwneg73_83 in73 sn83 11140.846016
Rwneg73_84 in73 sn84 11140.846016
Rwneg73_85 in73 sn85 3183.098862
Rwneg73_86 in73 sn86 11140.846016
Rwneg73_87 in73 sn87 11140.846016
Rwneg73_88 in73 sn88 11140.846016
Rwneg73_89 in73 sn89 3183.098862
Rwneg73_90 in73 sn90 11140.846016
Rwneg73_91 in73 sn91 11140.846016
Rwneg73_92 in73 sn92 3183.098862
Rwneg73_93 in73 sn93 11140.846016
Rwneg73_94 in73 sn94 11140.846016
Rwneg73_95 in73 sn95 3183.098862
Rwneg73_96 in73 sn96 3183.098862
Rwneg73_97 in73 sn97 11140.846016
Rwneg73_98 in73 sn98 3183.098862
Rwneg73_99 in73 sn99 11140.846016
Rwneg73_100 in73 sn100 11140.846016
Rwneg74_1 in74 sn1 11140.846016
Rwneg74_2 in74 sn2 11140.846016
Rwneg74_3 in74 sn3 11140.846016
Rwneg74_4 in74 sn4 3183.098862
Rwneg74_5 in74 sn5 11140.846016
Rwneg74_6 in74 sn6 3183.098862
Rwneg74_7 in74 sn7 11140.846016
Rwneg74_8 in74 sn8 3183.098862
Rwneg74_9 in74 sn9 11140.846016
Rwneg74_10 in74 sn10 11140.846016
Rwneg74_11 in74 sn11 11140.846016
Rwneg74_12 in74 sn12 3183.098862
Rwneg74_13 in74 sn13 11140.846016
Rwneg74_14 in74 sn14 3183.098862
Rwneg74_15 in74 sn15 3183.098862
Rwneg74_16 in74 sn16 11140.846016
Rwneg74_17 in74 sn17 11140.846016
Rwneg74_18 in74 sn18 3183.098862
Rwneg74_19 in74 sn19 11140.846016
Rwneg74_20 in74 sn20 11140.846016
Rwneg74_21 in74 sn21 3183.098862
Rwneg74_22 in74 sn22 11140.846016
Rwneg74_23 in74 sn23 11140.846016
Rwneg74_24 in74 sn24 3183.098862
Rwneg74_25 in74 sn25 11140.846016
Rwneg74_26 in74 sn26 11140.846016
Rwneg74_27 in74 sn27 3183.098862
Rwneg74_28 in74 sn28 3183.098862
Rwneg74_29 in74 sn29 11140.846016
Rwneg74_30 in74 sn30 3183.098862
Rwneg74_31 in74 sn31 3183.098862
Rwneg74_32 in74 sn32 11140.846016
Rwneg74_33 in74 sn33 11140.846016
Rwneg74_34 in74 sn34 11140.846016
Rwneg74_35 in74 sn35 11140.846016
Rwneg74_36 in74 sn36 3183.098862
Rwneg74_37 in74 sn37 11140.846016
Rwneg74_38 in74 sn38 11140.846016
Rwneg74_39 in74 sn39 11140.846016
Rwneg74_40 in74 sn40 3183.098862
Rwneg74_41 in74 sn41 11140.846016
Rwneg74_42 in74 sn42 11140.846016
Rwneg74_43 in74 sn43 11140.846016
Rwneg74_44 in74 sn44 3183.098862
Rwneg74_45 in74 sn45 11140.846016
Rwneg74_46 in74 sn46 3183.098862
Rwneg74_47 in74 sn47 3183.098862
Rwneg74_48 in74 sn48 11140.846016
Rwneg74_49 in74 sn49 11140.846016
Rwneg74_50 in74 sn50 3183.098862
Rwneg74_51 in74 sn51 3183.098862
Rwneg74_52 in74 sn52 3183.098862
Rwneg74_53 in74 sn53 11140.846016
Rwneg74_54 in74 sn54 11140.846016
Rwneg74_55 in74 sn55 11140.846016
Rwneg74_56 in74 sn56 11140.846016
Rwneg74_57 in74 sn57 3183.098862
Rwneg74_58 in74 sn58 3183.098862
Rwneg74_59 in74 sn59 11140.846016
Rwneg74_60 in74 sn60 3183.098862
Rwneg74_61 in74 sn61 11140.846016
Rwneg74_62 in74 sn62 3183.098862
Rwneg74_63 in74 sn63 3183.098862
Rwneg74_64 in74 sn64 3183.098862
Rwneg74_65 in74 sn65 11140.846016
Rwneg74_66 in74 sn66 11140.846016
Rwneg74_67 in74 sn67 11140.846016
Rwneg74_68 in74 sn68 11140.846016
Rwneg74_69 in74 sn69 11140.846016
Rwneg74_70 in74 sn70 3183.098862
Rwneg74_71 in74 sn71 3183.098862
Rwneg74_72 in74 sn72 11140.846016
Rwneg74_73 in74 sn73 11140.846016
Rwneg74_74 in74 sn74 3183.098862
Rwneg74_75 in74 sn75 11140.846016
Rwneg74_76 in74 sn76 3183.098862
Rwneg74_77 in74 sn77 11140.846016
Rwneg74_78 in74 sn78 3183.098862
Rwneg74_79 in74 sn79 11140.846016
Rwneg74_80 in74 sn80 3183.098862
Rwneg74_81 in74 sn81 11140.846016
Rwneg74_82 in74 sn82 11140.846016
Rwneg74_83 in74 sn83 3183.098862
Rwneg74_84 in74 sn84 11140.846016
Rwneg74_85 in74 sn85 11140.846016
Rwneg74_86 in74 sn86 11140.846016
Rwneg74_87 in74 sn87 11140.846016
Rwneg74_88 in74 sn88 11140.846016
Rwneg74_89 in74 sn89 11140.846016
Rwneg74_90 in74 sn90 3183.098862
Rwneg74_91 in74 sn91 11140.846016
Rwneg74_92 in74 sn92 11140.846016
Rwneg74_93 in74 sn93 11140.846016
Rwneg74_94 in74 sn94 3183.098862
Rwneg74_95 in74 sn95 11140.846016
Rwneg74_96 in74 sn96 3183.098862
Rwneg74_97 in74 sn97 3183.098862
Rwneg74_98 in74 sn98 11140.846016
Rwneg74_99 in74 sn99 3183.098862
Rwneg74_100 in74 sn100 3183.098862
Rwneg75_1 in75 sn1 11140.846016
Rwneg75_2 in75 sn2 3183.098862
Rwneg75_3 in75 sn3 11140.846016
Rwneg75_4 in75 sn4 11140.846016
Rwneg75_5 in75 sn5 11140.846016
Rwneg75_6 in75 sn6 3183.098862
Rwneg75_7 in75 sn7 11140.846016
Rwneg75_8 in75 sn8 3183.098862
Rwneg75_9 in75 sn9 3183.098862
Rwneg75_10 in75 sn10 3183.098862
Rwneg75_11 in75 sn11 11140.846016
Rwneg75_12 in75 sn12 11140.846016
Rwneg75_13 in75 sn13 3183.098862
Rwneg75_14 in75 sn14 11140.846016
Rwneg75_15 in75 sn15 11140.846016
Rwneg75_16 in75 sn16 3183.098862
Rwneg75_17 in75 sn17 11140.846016
Rwneg75_18 in75 sn18 3183.098862
Rwneg75_19 in75 sn19 11140.846016
Rwneg75_20 in75 sn20 11140.846016
Rwneg75_21 in75 sn21 3183.098862
Rwneg75_22 in75 sn22 11140.846016
Rwneg75_23 in75 sn23 11140.846016
Rwneg75_24 in75 sn24 11140.846016
Rwneg75_25 in75 sn25 3183.098862
Rwneg75_26 in75 sn26 3183.098862
Rwneg75_27 in75 sn27 11140.846016
Rwneg75_28 in75 sn28 3183.098862
Rwneg75_29 in75 sn29 3183.098862
Rwneg75_30 in75 sn30 11140.846016
Rwneg75_31 in75 sn31 11140.846016
Rwneg75_32 in75 sn32 3183.098862
Rwneg75_33 in75 sn33 11140.846016
Rwneg75_34 in75 sn34 11140.846016
Rwneg75_35 in75 sn35 3183.098862
Rwneg75_36 in75 sn36 11140.846016
Rwneg75_37 in75 sn37 11140.846016
Rwneg75_38 in75 sn38 11140.846016
Rwneg75_39 in75 sn39 11140.846016
Rwneg75_40 in75 sn40 3183.098862
Rwneg75_41 in75 sn41 3183.098862
Rwneg75_42 in75 sn42 11140.846016
Rwneg75_43 in75 sn43 11140.846016
Rwneg75_44 in75 sn44 3183.098862
Rwneg75_45 in75 sn45 11140.846016
Rwneg75_46 in75 sn46 11140.846016
Rwneg75_47 in75 sn47 3183.098862
Rwneg75_48 in75 sn48 3183.098862
Rwneg75_49 in75 sn49 11140.846016
Rwneg75_50 in75 sn50 11140.846016
Rwneg75_51 in75 sn51 11140.846016
Rwneg75_52 in75 sn52 11140.846016
Rwneg75_53 in75 sn53 11140.846016
Rwneg75_54 in75 sn54 11140.846016
Rwneg75_55 in75 sn55 11140.846016
Rwneg75_56 in75 sn56 11140.846016
Rwneg75_57 in75 sn57 3183.098862
Rwneg75_58 in75 sn58 3183.098862
Rwneg75_59 in75 sn59 11140.846016
Rwneg75_60 in75 sn60 11140.846016
Rwneg75_61 in75 sn61 3183.098862
Rwneg75_62 in75 sn62 3183.098862
Rwneg75_63 in75 sn63 11140.846016
Rwneg75_64 in75 sn64 3183.098862
Rwneg75_65 in75 sn65 11140.846016
Rwneg75_66 in75 sn66 3183.098862
Rwneg75_67 in75 sn67 3183.098862
Rwneg75_68 in75 sn68 11140.846016
Rwneg75_69 in75 sn69 11140.846016
Rwneg75_70 in75 sn70 11140.846016
Rwneg75_71 in75 sn71 3183.098862
Rwneg75_72 in75 sn72 11140.846016
Rwneg75_73 in75 sn73 3183.098862
Rwneg75_74 in75 sn74 11140.846016
Rwneg75_75 in75 sn75 11140.846016
Rwneg75_76 in75 sn76 3183.098862
Rwneg75_77 in75 sn77 11140.846016
Rwneg75_78 in75 sn78 3183.098862
Rwneg75_79 in75 sn79 11140.846016
Rwneg75_80 in75 sn80 11140.846016
Rwneg75_81 in75 sn81 3183.098862
Rwneg75_82 in75 sn82 3183.098862
Rwneg75_83 in75 sn83 11140.846016
Rwneg75_84 in75 sn84 11140.846016
Rwneg75_85 in75 sn85 11140.846016
Rwneg75_86 in75 sn86 11140.846016
Rwneg75_87 in75 sn87 3183.098862
Rwneg75_88 in75 sn88 11140.846016
Rwneg75_89 in75 sn89 3183.098862
Rwneg75_90 in75 sn90 3183.098862
Rwneg75_91 in75 sn91 11140.846016
Rwneg75_92 in75 sn92 11140.846016
Rwneg75_93 in75 sn93 11140.846016
Rwneg75_94 in75 sn94 3183.098862
Rwneg75_95 in75 sn95 11140.846016
Rwneg75_96 in75 sn96 3183.098862
Rwneg75_97 in75 sn97 3183.098862
Rwneg75_98 in75 sn98 3183.098862
Rwneg75_99 in75 sn99 11140.846016
Rwneg75_100 in75 sn100 3183.098862
Rwneg76_1 in76 sn1 11140.846016
Rwneg76_2 in76 sn2 11140.846016
Rwneg76_3 in76 sn3 3183.098862
Rwneg76_4 in76 sn4 3183.098862
Rwneg76_5 in76 sn5 3183.098862
Rwneg76_6 in76 sn6 11140.846016
Rwneg76_7 in76 sn7 11140.846016
Rwneg76_8 in76 sn8 3183.098862
Rwneg76_9 in76 sn9 11140.846016
Rwneg76_10 in76 sn10 3183.098862
Rwneg76_11 in76 sn11 11140.846016
Rwneg76_12 in76 sn12 3183.098862
Rwneg76_13 in76 sn13 11140.846016
Rwneg76_14 in76 sn14 11140.846016
Rwneg76_15 in76 sn15 3183.098862
Rwneg76_16 in76 sn16 3183.098862
Rwneg76_17 in76 sn17 11140.846016
Rwneg76_18 in76 sn18 11140.846016
Rwneg76_19 in76 sn19 3183.098862
Rwneg76_20 in76 sn20 3183.098862
Rwneg76_21 in76 sn21 3183.098862
Rwneg76_22 in76 sn22 3183.098862
Rwneg76_23 in76 sn23 11140.846016
Rwneg76_24 in76 sn24 11140.846016
Rwneg76_25 in76 sn25 11140.846016
Rwneg76_26 in76 sn26 3183.098862
Rwneg76_27 in76 sn27 3183.098862
Rwneg76_28 in76 sn28 11140.846016
Rwneg76_29 in76 sn29 3183.098862
Rwneg76_30 in76 sn30 3183.098862
Rwneg76_31 in76 sn31 11140.846016
Rwneg76_32 in76 sn32 11140.846016
Rwneg76_33 in76 sn33 11140.846016
Rwneg76_34 in76 sn34 11140.846016
Rwneg76_35 in76 sn35 3183.098862
Rwneg76_36 in76 sn36 3183.098862
Rwneg76_37 in76 sn37 11140.846016
Rwneg76_38 in76 sn38 11140.846016
Rwneg76_39 in76 sn39 11140.846016
Rwneg76_40 in76 sn40 11140.846016
Rwneg76_41 in76 sn41 3183.098862
Rwneg76_42 in76 sn42 3183.098862
Rwneg76_43 in76 sn43 11140.846016
Rwneg76_44 in76 sn44 3183.098862
Rwneg76_45 in76 sn45 3183.098862
Rwneg76_46 in76 sn46 11140.846016
Rwneg76_47 in76 sn47 11140.846016
Rwneg76_48 in76 sn48 3183.098862
Rwneg76_49 in76 sn49 11140.846016
Rwneg76_50 in76 sn50 11140.846016
Rwneg76_51 in76 sn51 3183.098862
Rwneg76_52 in76 sn52 11140.846016
Rwneg76_53 in76 sn53 11140.846016
Rwneg76_54 in76 sn54 3183.098862
Rwneg76_55 in76 sn55 3183.098862
Rwneg76_56 in76 sn56 3183.098862
Rwneg76_57 in76 sn57 11140.846016
Rwneg76_58 in76 sn58 3183.098862
Rwneg76_59 in76 sn59 11140.846016
Rwneg76_60 in76 sn60 3183.098862
Rwneg76_61 in76 sn61 3183.098862
Rwneg76_62 in76 sn62 11140.846016
Rwneg76_63 in76 sn63 3183.098862
Rwneg76_64 in76 sn64 3183.098862
Rwneg76_65 in76 sn65 11140.846016
Rwneg76_66 in76 sn66 3183.098862
Rwneg76_67 in76 sn67 11140.846016
Rwneg76_68 in76 sn68 3183.098862
Rwneg76_69 in76 sn69 11140.846016
Rwneg76_70 in76 sn70 11140.846016
Rwneg76_71 in76 sn71 11140.846016
Rwneg76_72 in76 sn72 11140.846016
Rwneg76_73 in76 sn73 3183.098862
Rwneg76_74 in76 sn74 11140.846016
Rwneg76_75 in76 sn75 11140.846016
Rwneg76_76 in76 sn76 11140.846016
Rwneg76_77 in76 sn77 11140.846016
Rwneg76_78 in76 sn78 11140.846016
Rwneg76_79 in76 sn79 3183.098862
Rwneg76_80 in76 sn80 11140.846016
Rwneg76_81 in76 sn81 3183.098862
Rwneg76_82 in76 sn82 3183.098862
Rwneg76_83 in76 sn83 11140.846016
Rwneg76_84 in76 sn84 3183.098862
Rwneg76_85 in76 sn85 11140.846016
Rwneg76_86 in76 sn86 11140.846016
Rwneg76_87 in76 sn87 3183.098862
Rwneg76_88 in76 sn88 11140.846016
Rwneg76_89 in76 sn89 11140.846016
Rwneg76_90 in76 sn90 11140.846016
Rwneg76_91 in76 sn91 11140.846016
Rwneg76_92 in76 sn92 11140.846016
Rwneg76_93 in76 sn93 3183.098862
Rwneg76_94 in76 sn94 3183.098862
Rwneg76_95 in76 sn95 11140.846016
Rwneg76_96 in76 sn96 3183.098862
Rwneg76_97 in76 sn97 11140.846016
Rwneg76_98 in76 sn98 3183.098862
Rwneg76_99 in76 sn99 11140.846016
Rwneg76_100 in76 sn100 11140.846016
Rwneg77_1 in77 sn1 3183.098862
Rwneg77_2 in77 sn2 11140.846016
Rwneg77_3 in77 sn3 3183.098862
Rwneg77_4 in77 sn4 11140.846016
Rwneg77_5 in77 sn5 11140.846016
Rwneg77_6 in77 sn6 3183.098862
Rwneg77_7 in77 sn7 3183.098862
Rwneg77_8 in77 sn8 3183.098862
Rwneg77_9 in77 sn9 11140.846016
Rwneg77_10 in77 sn10 11140.846016
Rwneg77_11 in77 sn11 3183.098862
Rwneg77_12 in77 sn12 11140.846016
Rwneg77_13 in77 sn13 11140.846016
Rwneg77_14 in77 sn14 11140.846016
Rwneg77_15 in77 sn15 3183.098862
Rwneg77_16 in77 sn16 11140.846016
Rwneg77_17 in77 sn17 11140.846016
Rwneg77_18 in77 sn18 3183.098862
Rwneg77_19 in77 sn19 11140.846016
Rwneg77_20 in77 sn20 3183.098862
Rwneg77_21 in77 sn21 3183.098862
Rwneg77_22 in77 sn22 3183.098862
Rwneg77_23 in77 sn23 3183.098862
Rwneg77_24 in77 sn24 3183.098862
Rwneg77_25 in77 sn25 11140.846016
Rwneg77_26 in77 sn26 3183.098862
Rwneg77_27 in77 sn27 11140.846016
Rwneg77_28 in77 sn28 3183.098862
Rwneg77_29 in77 sn29 11140.846016
Rwneg77_30 in77 sn30 3183.098862
Rwneg77_31 in77 sn31 11140.846016
Rwneg77_32 in77 sn32 3183.098862
Rwneg77_33 in77 sn33 3183.098862
Rwneg77_34 in77 sn34 11140.846016
Rwneg77_35 in77 sn35 11140.846016
Rwneg77_36 in77 sn36 3183.098862
Rwneg77_37 in77 sn37 3183.098862
Rwneg77_38 in77 sn38 3183.098862
Rwneg77_39 in77 sn39 11140.846016
Rwneg77_40 in77 sn40 11140.846016
Rwneg77_41 in77 sn41 3183.098862
Rwneg77_42 in77 sn42 11140.846016
Rwneg77_43 in77 sn43 3183.098862
Rwneg77_44 in77 sn44 3183.098862
Rwneg77_45 in77 sn45 3183.098862
Rwneg77_46 in77 sn46 11140.846016
Rwneg77_47 in77 sn47 3183.098862
Rwneg77_48 in77 sn48 11140.846016
Rwneg77_49 in77 sn49 11140.846016
Rwneg77_50 in77 sn50 11140.846016
Rwneg77_51 in77 sn51 11140.846016
Rwneg77_52 in77 sn52 11140.846016
Rwneg77_53 in77 sn53 3183.098862
Rwneg77_54 in77 sn54 11140.846016
Rwneg77_55 in77 sn55 11140.846016
Rwneg77_56 in77 sn56 11140.846016
Rwneg77_57 in77 sn57 11140.846016
Rwneg77_58 in77 sn58 11140.846016
Rwneg77_59 in77 sn59 3183.098862
Rwneg77_60 in77 sn60 11140.846016
Rwneg77_61 in77 sn61 3183.098862
Rwneg77_62 in77 sn62 11140.846016
Rwneg77_63 in77 sn63 11140.846016
Rwneg77_64 in77 sn64 3183.098862
Rwneg77_65 in77 sn65 11140.846016
Rwneg77_66 in77 sn66 11140.846016
Rwneg77_67 in77 sn67 3183.098862
Rwneg77_68 in77 sn68 3183.098862
Rwneg77_69 in77 sn69 11140.846016
Rwneg77_70 in77 sn70 3183.098862
Rwneg77_71 in77 sn71 11140.846016
Rwneg77_72 in77 sn72 11140.846016
Rwneg77_73 in77 sn73 11140.846016
Rwneg77_74 in77 sn74 3183.098862
Rwneg77_75 in77 sn75 3183.098862
Rwneg77_76 in77 sn76 3183.098862
Rwneg77_77 in77 sn77 11140.846016
Rwneg77_78 in77 sn78 11140.846016
Rwneg77_79 in77 sn79 11140.846016
Rwneg77_80 in77 sn80 11140.846016
Rwneg77_81 in77 sn81 3183.098862
Rwneg77_82 in77 sn82 11140.846016
Rwneg77_83 in77 sn83 11140.846016
Rwneg77_84 in77 sn84 11140.846016
Rwneg77_85 in77 sn85 11140.846016
Rwneg77_86 in77 sn86 11140.846016
Rwneg77_87 in77 sn87 11140.846016
Rwneg77_88 in77 sn88 11140.846016
Rwneg77_89 in77 sn89 3183.098862
Rwneg77_90 in77 sn90 3183.098862
Rwneg77_91 in77 sn91 3183.098862
Rwneg77_92 in77 sn92 3183.098862
Rwneg77_93 in77 sn93 11140.846016
Rwneg77_94 in77 sn94 3183.098862
Rwneg77_95 in77 sn95 11140.846016
Rwneg77_96 in77 sn96 3183.098862
Rwneg77_97 in77 sn97 3183.098862
Rwneg77_98 in77 sn98 11140.846016
Rwneg77_99 in77 sn99 11140.846016
Rwneg77_100 in77 sn100 3183.098862
Rwneg78_1 in78 sn1 11140.846016
Rwneg78_2 in78 sn2 11140.846016
Rwneg78_3 in78 sn3 11140.846016
Rwneg78_4 in78 sn4 11140.846016
Rwneg78_5 in78 sn5 3183.098862
Rwneg78_6 in78 sn6 11140.846016
Rwneg78_7 in78 sn7 3183.098862
Rwneg78_8 in78 sn8 3183.098862
Rwneg78_9 in78 sn9 11140.846016
Rwneg78_10 in78 sn10 11140.846016
Rwneg78_11 in78 sn11 3183.098862
Rwneg78_12 in78 sn12 3183.098862
Rwneg78_13 in78 sn13 11140.846016
Rwneg78_14 in78 sn14 11140.846016
Rwneg78_15 in78 sn15 11140.846016
Rwneg78_16 in78 sn16 11140.846016
Rwneg78_17 in78 sn17 11140.846016
Rwneg78_18 in78 sn18 11140.846016
Rwneg78_19 in78 sn19 3183.098862
Rwneg78_20 in78 sn20 3183.098862
Rwneg78_21 in78 sn21 3183.098862
Rwneg78_22 in78 sn22 3183.098862
Rwneg78_23 in78 sn23 3183.098862
Rwneg78_24 in78 sn24 3183.098862
Rwneg78_25 in78 sn25 11140.846016
Rwneg78_26 in78 sn26 11140.846016
Rwneg78_27 in78 sn27 3183.098862
Rwneg78_28 in78 sn28 3183.098862
Rwneg78_29 in78 sn29 11140.846016
Rwneg78_30 in78 sn30 3183.098862
Rwneg78_31 in78 sn31 3183.098862
Rwneg78_32 in78 sn32 11140.846016
Rwneg78_33 in78 sn33 11140.846016
Rwneg78_34 in78 sn34 11140.846016
Rwneg78_35 in78 sn35 3183.098862
Rwneg78_36 in78 sn36 3183.098862
Rwneg78_37 in78 sn37 11140.846016
Rwneg78_38 in78 sn38 3183.098862
Rwneg78_39 in78 sn39 3183.098862
Rwneg78_40 in78 sn40 3183.098862
Rwneg78_41 in78 sn41 11140.846016
Rwneg78_42 in78 sn42 11140.846016
Rwneg78_43 in78 sn43 3183.098862
Rwneg78_44 in78 sn44 11140.846016
Rwneg78_45 in78 sn45 11140.846016
Rwneg78_46 in78 sn46 11140.846016
Rwneg78_47 in78 sn47 3183.098862
Rwneg78_48 in78 sn48 11140.846016
Rwneg78_49 in78 sn49 3183.098862
Rwneg78_50 in78 sn50 11140.846016
Rwneg78_51 in78 sn51 11140.846016
Rwneg78_52 in78 sn52 3183.098862
Rwneg78_53 in78 sn53 3183.098862
Rwneg78_54 in78 sn54 3183.098862
Rwneg78_55 in78 sn55 11140.846016
Rwneg78_56 in78 sn56 11140.846016
Rwneg78_57 in78 sn57 11140.846016
Rwneg78_58 in78 sn58 11140.846016
Rwneg78_59 in78 sn59 3183.098862
Rwneg78_60 in78 sn60 3183.098862
Rwneg78_61 in78 sn61 11140.846016
Rwneg78_62 in78 sn62 3183.098862
Rwneg78_63 in78 sn63 3183.098862
Rwneg78_64 in78 sn64 11140.846016
Rwneg78_65 in78 sn65 11140.846016
Rwneg78_66 in78 sn66 11140.846016
Rwneg78_67 in78 sn67 11140.846016
Rwneg78_68 in78 sn68 3183.098862
Rwneg78_69 in78 sn69 11140.846016
Rwneg78_70 in78 sn70 3183.098862
Rwneg78_71 in78 sn71 11140.846016
Rwneg78_72 in78 sn72 11140.846016
Rwneg78_73 in78 sn73 11140.846016
Rwneg78_74 in78 sn74 3183.098862
Rwneg78_75 in78 sn75 3183.098862
Rwneg78_76 in78 sn76 3183.098862
Rwneg78_77 in78 sn77 11140.846016
Rwneg78_78 in78 sn78 3183.098862
Rwneg78_79 in78 sn79 3183.098862
Rwneg78_80 in78 sn80 11140.846016
Rwneg78_81 in78 sn81 11140.846016
Rwneg78_82 in78 sn82 11140.846016
Rwneg78_83 in78 sn83 11140.846016
Rwneg78_84 in78 sn84 11140.846016
Rwneg78_85 in78 sn85 11140.846016
Rwneg78_86 in78 sn86 11140.846016
Rwneg78_87 in78 sn87 11140.846016
Rwneg78_88 in78 sn88 3183.098862
Rwneg78_89 in78 sn89 11140.846016
Rwneg78_90 in78 sn90 3183.098862
Rwneg78_91 in78 sn91 11140.846016
Rwneg78_92 in78 sn92 3183.098862
Rwneg78_93 in78 sn93 11140.846016
Rwneg78_94 in78 sn94 3183.098862
Rwneg78_95 in78 sn95 3183.098862
Rwneg78_96 in78 sn96 11140.846016
Rwneg78_97 in78 sn97 11140.846016
Rwneg78_98 in78 sn98 11140.846016
Rwneg78_99 in78 sn99 11140.846016
Rwneg78_100 in78 sn100 3183.098862
Rwneg79_1 in79 sn1 11140.846016
Rwneg79_2 in79 sn2 3183.098862
Rwneg79_3 in79 sn3 11140.846016
Rwneg79_4 in79 sn4 3183.098862
Rwneg79_5 in79 sn5 3183.098862
Rwneg79_6 in79 sn6 3183.098862
Rwneg79_7 in79 sn7 11140.846016
Rwneg79_8 in79 sn8 3183.098862
Rwneg79_9 in79 sn9 11140.846016
Rwneg79_10 in79 sn10 3183.098862
Rwneg79_11 in79 sn11 3183.098862
Rwneg79_12 in79 sn12 3183.098862
Rwneg79_13 in79 sn13 3183.098862
Rwneg79_14 in79 sn14 11140.846016
Rwneg79_15 in79 sn15 11140.846016
Rwneg79_16 in79 sn16 11140.846016
Rwneg79_17 in79 sn17 11140.846016
Rwneg79_18 in79 sn18 3183.098862
Rwneg79_19 in79 sn19 11140.846016
Rwneg79_20 in79 sn20 11140.846016
Rwneg79_21 in79 sn21 3183.098862
Rwneg79_22 in79 sn22 3183.098862
Rwneg79_23 in79 sn23 11140.846016
Rwneg79_24 in79 sn24 3183.098862
Rwneg79_25 in79 sn25 11140.846016
Rwneg79_26 in79 sn26 3183.098862
Rwneg79_27 in79 sn27 11140.846016
Rwneg79_28 in79 sn28 3183.098862
Rwneg79_29 in79 sn29 3183.098862
Rwneg79_30 in79 sn30 11140.846016
Rwneg79_31 in79 sn31 3183.098862
Rwneg79_32 in79 sn32 3183.098862
Rwneg79_33 in79 sn33 11140.846016
Rwneg79_34 in79 sn34 3183.098862
Rwneg79_35 in79 sn35 3183.098862
Rwneg79_36 in79 sn36 11140.846016
Rwneg79_37 in79 sn37 3183.098862
Rwneg79_38 in79 sn38 3183.098862
Rwneg79_39 in79 sn39 11140.846016
Rwneg79_40 in79 sn40 3183.098862
Rwneg79_41 in79 sn41 11140.846016
Rwneg79_42 in79 sn42 3183.098862
Rwneg79_43 in79 sn43 11140.846016
Rwneg79_44 in79 sn44 3183.098862
Rwneg79_45 in79 sn45 3183.098862
Rwneg79_46 in79 sn46 11140.846016
Rwneg79_47 in79 sn47 3183.098862
Rwneg79_48 in79 sn48 3183.098862
Rwneg79_49 in79 sn49 11140.846016
Rwneg79_50 in79 sn50 3183.098862
Rwneg79_51 in79 sn51 3183.098862
Rwneg79_52 in79 sn52 11140.846016
Rwneg79_53 in79 sn53 11140.846016
Rwneg79_54 in79 sn54 3183.098862
Rwneg79_55 in79 sn55 11140.846016
Rwneg79_56 in79 sn56 3183.098862
Rwneg79_57 in79 sn57 11140.846016
Rwneg79_58 in79 sn58 11140.846016
Rwneg79_59 in79 sn59 11140.846016
Rwneg79_60 in79 sn60 3183.098862
Rwneg79_61 in79 sn61 3183.098862
Rwneg79_62 in79 sn62 11140.846016
Rwneg79_63 in79 sn63 11140.846016
Rwneg79_64 in79 sn64 3183.098862
Rwneg79_65 in79 sn65 11140.846016
Rwneg79_66 in79 sn66 3183.098862
Rwneg79_67 in79 sn67 3183.098862
Rwneg79_68 in79 sn68 3183.098862
Rwneg79_69 in79 sn69 11140.846016
Rwneg79_70 in79 sn70 11140.846016
Rwneg79_71 in79 sn71 11140.846016
Rwneg79_72 in79 sn72 3183.098862
Rwneg79_73 in79 sn73 3183.098862
Rwneg79_74 in79 sn74 11140.846016
Rwneg79_75 in79 sn75 3183.098862
Rwneg79_76 in79 sn76 11140.846016
Rwneg79_77 in79 sn77 3183.098862
Rwneg79_78 in79 sn78 11140.846016
Rwneg79_79 in79 sn79 11140.846016
Rwneg79_80 in79 sn80 3183.098862
Rwneg79_81 in79 sn81 11140.846016
Rwneg79_82 in79 sn82 3183.098862
Rwneg79_83 in79 sn83 3183.098862
Rwneg79_84 in79 sn84 11140.846016
Rwneg79_85 in79 sn85 3183.098862
Rwneg79_86 in79 sn86 11140.846016
Rwneg79_87 in79 sn87 11140.846016
Rwneg79_88 in79 sn88 11140.846016
Rwneg79_89 in79 sn89 3183.098862
Rwneg79_90 in79 sn90 3183.098862
Rwneg79_91 in79 sn91 3183.098862
Rwneg79_92 in79 sn92 3183.098862
Rwneg79_93 in79 sn93 3183.098862
Rwneg79_94 in79 sn94 11140.846016
Rwneg79_95 in79 sn95 11140.846016
Rwneg79_96 in79 sn96 3183.098862
Rwneg79_97 in79 sn97 11140.846016
Rwneg79_98 in79 sn98 11140.846016
Rwneg79_99 in79 sn99 3183.098862
Rwneg79_100 in79 sn100 3183.098862
Rwneg80_1 in80 sn1 11140.846016
Rwneg80_2 in80 sn2 11140.846016
Rwneg80_3 in80 sn3 3183.098862
Rwneg80_4 in80 sn4 3183.098862
Rwneg80_5 in80 sn5 3183.098862
Rwneg80_6 in80 sn6 11140.846016
Rwneg80_7 in80 sn7 11140.846016
Rwneg80_8 in80 sn8 11140.846016
Rwneg80_9 in80 sn9 3183.098862
Rwneg80_10 in80 sn10 3183.098862
Rwneg80_11 in80 sn11 3183.098862
Rwneg80_12 in80 sn12 11140.846016
Rwneg80_13 in80 sn13 3183.098862
Rwneg80_14 in80 sn14 3183.098862
Rwneg80_15 in80 sn15 3183.098862
Rwneg80_16 in80 sn16 3183.098862
Rwneg80_17 in80 sn17 3183.098862
Rwneg80_18 in80 sn18 11140.846016
Rwneg80_19 in80 sn19 11140.846016
Rwneg80_20 in80 sn20 11140.846016
Rwneg80_21 in80 sn21 3183.098862
Rwneg80_22 in80 sn22 11140.846016
Rwneg80_23 in80 sn23 11140.846016
Rwneg80_24 in80 sn24 11140.846016
Rwneg80_25 in80 sn25 3183.098862
Rwneg80_26 in80 sn26 3183.098862
Rwneg80_27 in80 sn27 11140.846016
Rwneg80_28 in80 sn28 3183.098862
Rwneg80_29 in80 sn29 3183.098862
Rwneg80_30 in80 sn30 11140.846016
Rwneg80_31 in80 sn31 3183.098862
Rwneg80_32 in80 sn32 11140.846016
Rwneg80_33 in80 sn33 3183.098862
Rwneg80_34 in80 sn34 11140.846016
Rwneg80_35 in80 sn35 3183.098862
Rwneg80_36 in80 sn36 3183.098862
Rwneg80_37 in80 sn37 3183.098862
Rwneg80_38 in80 sn38 11140.846016
Rwneg80_39 in80 sn39 11140.846016
Rwneg80_40 in80 sn40 3183.098862
Rwneg80_41 in80 sn41 11140.846016
Rwneg80_42 in80 sn42 3183.098862
Rwneg80_43 in80 sn43 11140.846016
Rwneg80_44 in80 sn44 11140.846016
Rwneg80_45 in80 sn45 11140.846016
Rwneg80_46 in80 sn46 3183.098862
Rwneg80_47 in80 sn47 3183.098862
Rwneg80_48 in80 sn48 11140.846016
Rwneg80_49 in80 sn49 11140.846016
Rwneg80_50 in80 sn50 11140.846016
Rwneg80_51 in80 sn51 11140.846016
Rwneg80_52 in80 sn52 3183.098862
Rwneg80_53 in80 sn53 3183.098862
Rwneg80_54 in80 sn54 11140.846016
Rwneg80_55 in80 sn55 11140.846016
Rwneg80_56 in80 sn56 11140.846016
Rwneg80_57 in80 sn57 3183.098862
Rwneg80_58 in80 sn58 3183.098862
Rwneg80_59 in80 sn59 11140.846016
Rwneg80_60 in80 sn60 11140.846016
Rwneg80_61 in80 sn61 3183.098862
Rwneg80_62 in80 sn62 3183.098862
Rwneg80_63 in80 sn63 3183.098862
Rwneg80_64 in80 sn64 11140.846016
Rwneg80_65 in80 sn65 11140.846016
Rwneg80_66 in80 sn66 11140.846016
Rwneg80_67 in80 sn67 11140.846016
Rwneg80_68 in80 sn68 3183.098862
Rwneg80_69 in80 sn69 3183.098862
Rwneg80_70 in80 sn70 11140.846016
Rwneg80_71 in80 sn71 11140.846016
Rwneg80_72 in80 sn72 11140.846016
Rwneg80_73 in80 sn73 3183.098862
Rwneg80_74 in80 sn74 3183.098862
Rwneg80_75 in80 sn75 11140.846016
Rwneg80_76 in80 sn76 11140.846016
Rwneg80_77 in80 sn77 3183.098862
Rwneg80_78 in80 sn78 3183.098862
Rwneg80_79 in80 sn79 3183.098862
Rwneg80_80 in80 sn80 3183.098862
Rwneg80_81 in80 sn81 11140.846016
Rwneg80_82 in80 sn82 11140.846016
Rwneg80_83 in80 sn83 3183.098862
Rwneg80_84 in80 sn84 11140.846016
Rwneg80_85 in80 sn85 11140.846016
Rwneg80_86 in80 sn86 11140.846016
Rwneg80_87 in80 sn87 11140.846016
Rwneg80_88 in80 sn88 11140.846016
Rwneg80_89 in80 sn89 11140.846016
Rwneg80_90 in80 sn90 11140.846016
Rwneg80_91 in80 sn91 3183.098862
Rwneg80_92 in80 sn92 11140.846016
Rwneg80_93 in80 sn93 11140.846016
Rwneg80_94 in80 sn94 3183.098862
Rwneg80_95 in80 sn95 11140.846016
Rwneg80_96 in80 sn96 11140.846016
Rwneg80_97 in80 sn97 11140.846016
Rwneg80_98 in80 sn98 11140.846016
Rwneg80_99 in80 sn99 3183.098862
Rwneg80_100 in80 sn100 3183.098862
Rwneg81_1 in81 sn1 11140.846016
Rwneg81_2 in81 sn2 3183.098862
Rwneg81_3 in81 sn3 3183.098862
Rwneg81_4 in81 sn4 11140.846016
Rwneg81_5 in81 sn5 3183.098862
Rwneg81_6 in81 sn6 3183.098862
Rwneg81_7 in81 sn7 11140.846016
Rwneg81_8 in81 sn8 11140.846016
Rwneg81_9 in81 sn9 3183.098862
Rwneg81_10 in81 sn10 11140.846016
Rwneg81_11 in81 sn11 3183.098862
Rwneg81_12 in81 sn12 11140.846016
Rwneg81_13 in81 sn13 3183.098862
Rwneg81_14 in81 sn14 3183.098862
Rwneg81_15 in81 sn15 3183.098862
Rwneg81_16 in81 sn16 11140.846016
Rwneg81_17 in81 sn17 11140.846016
Rwneg81_18 in81 sn18 11140.846016
Rwneg81_19 in81 sn19 11140.846016
Rwneg81_20 in81 sn20 11140.846016
Rwneg81_21 in81 sn21 3183.098862
Rwneg81_22 in81 sn22 11140.846016
Rwneg81_23 in81 sn23 3183.098862
Rwneg81_24 in81 sn24 11140.846016
Rwneg81_25 in81 sn25 11140.846016
Rwneg81_26 in81 sn26 11140.846016
Rwneg81_27 in81 sn27 3183.098862
Rwneg81_28 in81 sn28 11140.846016
Rwneg81_29 in81 sn29 11140.846016
Rwneg81_30 in81 sn30 11140.846016
Rwneg81_31 in81 sn31 3183.098862
Rwneg81_32 in81 sn32 3183.098862
Rwneg81_33 in81 sn33 3183.098862
Rwneg81_34 in81 sn34 3183.098862
Rwneg81_35 in81 sn35 3183.098862
Rwneg81_36 in81 sn36 11140.846016
Rwneg81_37 in81 sn37 3183.098862
Rwneg81_38 in81 sn38 3183.098862
Rwneg81_39 in81 sn39 3183.098862
Rwneg81_40 in81 sn40 11140.846016
Rwneg81_41 in81 sn41 11140.846016
Rwneg81_42 in81 sn42 11140.846016
Rwneg81_43 in81 sn43 11140.846016
Rwneg81_44 in81 sn44 3183.098862
Rwneg81_45 in81 sn45 11140.846016
Rwneg81_46 in81 sn46 3183.098862
Rwneg81_47 in81 sn47 3183.098862
Rwneg81_48 in81 sn48 3183.098862
Rwneg81_49 in81 sn49 11140.846016
Rwneg81_50 in81 sn50 3183.098862
Rwneg81_51 in81 sn51 11140.846016
Rwneg81_52 in81 sn52 11140.846016
Rwneg81_53 in81 sn53 3183.098862
Rwneg81_54 in81 sn54 11140.846016
Rwneg81_55 in81 sn55 3183.098862
Rwneg81_56 in81 sn56 3183.098862
Rwneg81_57 in81 sn57 3183.098862
Rwneg81_58 in81 sn58 3183.098862
Rwneg81_59 in81 sn59 11140.846016
Rwneg81_60 in81 sn60 3183.098862
Rwneg81_61 in81 sn61 3183.098862
Rwneg81_62 in81 sn62 3183.098862
Rwneg81_63 in81 sn63 11140.846016
Rwneg81_64 in81 sn64 3183.098862
Rwneg81_65 in81 sn65 11140.846016
Rwneg81_66 in81 sn66 11140.846016
Rwneg81_67 in81 sn67 11140.846016
Rwneg81_68 in81 sn68 11140.846016
Rwneg81_69 in81 sn69 11140.846016
Rwneg81_70 in81 sn70 11140.846016
Rwneg81_71 in81 sn71 3183.098862
Rwneg81_72 in81 sn72 11140.846016
Rwneg81_73 in81 sn73 11140.846016
Rwneg81_74 in81 sn74 3183.098862
Rwneg81_75 in81 sn75 11140.846016
Rwneg81_76 in81 sn76 11140.846016
Rwneg81_77 in81 sn77 3183.098862
Rwneg81_78 in81 sn78 3183.098862
Rwneg81_79 in81 sn79 3183.098862
Rwneg81_80 in81 sn80 3183.098862
Rwneg81_81 in81 sn81 11140.846016
Rwneg81_82 in81 sn82 3183.098862
Rwneg81_83 in81 sn83 11140.846016
Rwneg81_84 in81 sn84 11140.846016
Rwneg81_85 in81 sn85 11140.846016
Rwneg81_86 in81 sn86 11140.846016
Rwneg81_87 in81 sn87 11140.846016
Rwneg81_88 in81 sn88 3183.098862
Rwneg81_89 in81 sn89 3183.098862
Rwneg81_90 in81 sn90 11140.846016
Rwneg81_91 in81 sn91 11140.846016
Rwneg81_92 in81 sn92 3183.098862
Rwneg81_93 in81 sn93 3183.098862
Rwneg81_94 in81 sn94 3183.098862
Rwneg81_95 in81 sn95 11140.846016
Rwneg81_96 in81 sn96 3183.098862
Rwneg81_97 in81 sn97 3183.098862
Rwneg81_98 in81 sn98 3183.098862
Rwneg81_99 in81 sn99 3183.098862
Rwneg81_100 in81 sn100 3183.098862
Rwneg82_1 in82 sn1 3183.098862
Rwneg82_2 in82 sn2 11140.846016
Rwneg82_3 in82 sn3 3183.098862
Rwneg82_4 in82 sn4 11140.846016
Rwneg82_5 in82 sn5 3183.098862
Rwneg82_6 in82 sn6 3183.098862
Rwneg82_7 in82 sn7 11140.846016
Rwneg82_8 in82 sn8 11140.846016
Rwneg82_9 in82 sn9 11140.846016
Rwneg82_10 in82 sn10 11140.846016
Rwneg82_11 in82 sn11 3183.098862
Rwneg82_12 in82 sn12 3183.098862
Rwneg82_13 in82 sn13 3183.098862
Rwneg82_14 in82 sn14 11140.846016
Rwneg82_15 in82 sn15 3183.098862
Rwneg82_16 in82 sn16 11140.846016
Rwneg82_17 in82 sn17 3183.098862
Rwneg82_18 in82 sn18 3183.098862
Rwneg82_19 in82 sn19 11140.846016
Rwneg82_20 in82 sn20 3183.098862
Rwneg82_21 in82 sn21 3183.098862
Rwneg82_22 in82 sn22 3183.098862
Rwneg82_23 in82 sn23 11140.846016
Rwneg82_24 in82 sn24 11140.846016
Rwneg82_25 in82 sn25 11140.846016
Rwneg82_26 in82 sn26 11140.846016
Rwneg82_27 in82 sn27 11140.846016
Rwneg82_28 in82 sn28 3183.098862
Rwneg82_29 in82 sn29 3183.098862
Rwneg82_30 in82 sn30 11140.846016
Rwneg82_31 in82 sn31 3183.098862
Rwneg82_32 in82 sn32 3183.098862
Rwneg82_33 in82 sn33 3183.098862
Rwneg82_34 in82 sn34 3183.098862
Rwneg82_35 in82 sn35 11140.846016
Rwneg82_36 in82 sn36 3183.098862
Rwneg82_37 in82 sn37 11140.846016
Rwneg82_38 in82 sn38 11140.846016
Rwneg82_39 in82 sn39 3183.098862
Rwneg82_40 in82 sn40 3183.098862
Rwneg82_41 in82 sn41 3183.098862
Rwneg82_42 in82 sn42 3183.098862
Rwneg82_43 in82 sn43 3183.098862
Rwneg82_44 in82 sn44 11140.846016
Rwneg82_45 in82 sn45 11140.846016
Rwneg82_46 in82 sn46 3183.098862
Rwneg82_47 in82 sn47 11140.846016
Rwneg82_48 in82 sn48 11140.846016
Rwneg82_49 in82 sn49 11140.846016
Rwneg82_50 in82 sn50 11140.846016
Rwneg82_51 in82 sn51 11140.846016
Rwneg82_52 in82 sn52 3183.098862
Rwneg82_53 in82 sn53 11140.846016
Rwneg82_54 in82 sn54 11140.846016
Rwneg82_55 in82 sn55 3183.098862
Rwneg82_56 in82 sn56 3183.098862
Rwneg82_57 in82 sn57 11140.846016
Rwneg82_58 in82 sn58 11140.846016
Rwneg82_59 in82 sn59 3183.098862
Rwneg82_60 in82 sn60 3183.098862
Rwneg82_61 in82 sn61 11140.846016
Rwneg82_62 in82 sn62 11140.846016
Rwneg82_63 in82 sn63 11140.846016
Rwneg82_64 in82 sn64 11140.846016
Rwneg82_65 in82 sn65 11140.846016
Rwneg82_66 in82 sn66 3183.098862
Rwneg82_67 in82 sn67 3183.098862
Rwneg82_68 in82 sn68 11140.846016
Rwneg82_69 in82 sn69 3183.098862
Rwneg82_70 in82 sn70 11140.846016
Rwneg82_71 in82 sn71 3183.098862
Rwneg82_72 in82 sn72 3183.098862
Rwneg82_73 in82 sn73 3183.098862
Rwneg82_74 in82 sn74 11140.846016
Rwneg82_75 in82 sn75 3183.098862
Rwneg82_76 in82 sn76 3183.098862
Rwneg82_77 in82 sn77 11140.846016
Rwneg82_78 in82 sn78 3183.098862
Rwneg82_79 in82 sn79 11140.846016
Rwneg82_80 in82 sn80 11140.846016
Rwneg82_81 in82 sn81 11140.846016
Rwneg82_82 in82 sn82 3183.098862
Rwneg82_83 in82 sn83 11140.846016
Rwneg82_84 in82 sn84 11140.846016
Rwneg82_85 in82 sn85 3183.098862
Rwneg82_86 in82 sn86 11140.846016
Rwneg82_87 in82 sn87 11140.846016
Rwneg82_88 in82 sn88 3183.098862
Rwneg82_89 in82 sn89 11140.846016
Rwneg82_90 in82 sn90 3183.098862
Rwneg82_91 in82 sn91 3183.098862
Rwneg82_92 in82 sn92 3183.098862
Rwneg82_93 in82 sn93 11140.846016
Rwneg82_94 in82 sn94 3183.098862
Rwneg82_95 in82 sn95 11140.846016
Rwneg82_96 in82 sn96 11140.846016
Rwneg82_97 in82 sn97 11140.846016
Rwneg82_98 in82 sn98 11140.846016
Rwneg82_99 in82 sn99 11140.846016
Rwneg82_100 in82 sn100 11140.846016
Rwneg83_1 in83 sn1 11140.846016
Rwneg83_2 in83 sn2 3183.098862
Rwneg83_3 in83 sn3 3183.098862
Rwneg83_4 in83 sn4 3183.098862
Rwneg83_5 in83 sn5 11140.846016
Rwneg83_6 in83 sn6 3183.098862
Rwneg83_7 in83 sn7 3183.098862
Rwneg83_8 in83 sn8 3183.098862
Rwneg83_9 in83 sn9 11140.846016
Rwneg83_10 in83 sn10 3183.098862
Rwneg83_11 in83 sn11 3183.098862
Rwneg83_12 in83 sn12 3183.098862
Rwneg83_13 in83 sn13 3183.098862
Rwneg83_14 in83 sn14 11140.846016
Rwneg83_15 in83 sn15 11140.846016
Rwneg83_16 in83 sn16 11140.846016
Rwneg83_17 in83 sn17 11140.846016
Rwneg83_18 in83 sn18 3183.098862
Rwneg83_19 in83 sn19 11140.846016
Rwneg83_20 in83 sn20 3183.098862
Rwneg83_21 in83 sn21 3183.098862
Rwneg83_22 in83 sn22 3183.098862
Rwneg83_23 in83 sn23 3183.098862
Rwneg83_24 in83 sn24 3183.098862
Rwneg83_25 in83 sn25 11140.846016
Rwneg83_26 in83 sn26 3183.098862
Rwneg83_27 in83 sn27 3183.098862
Rwneg83_28 in83 sn28 3183.098862
Rwneg83_29 in83 sn29 11140.846016
Rwneg83_30 in83 sn30 3183.098862
Rwneg83_31 in83 sn31 11140.846016
Rwneg83_32 in83 sn32 11140.846016
Rwneg83_33 in83 sn33 11140.846016
Rwneg83_34 in83 sn34 3183.098862
Rwneg83_35 in83 sn35 11140.846016
Rwneg83_36 in83 sn36 3183.098862
Rwneg83_37 in83 sn37 11140.846016
Rwneg83_38 in83 sn38 3183.098862
Rwneg83_39 in83 sn39 3183.098862
Rwneg83_40 in83 sn40 3183.098862
Rwneg83_41 in83 sn41 11140.846016
Rwneg83_42 in83 sn42 3183.098862
Rwneg83_43 in83 sn43 11140.846016
Rwneg83_44 in83 sn44 3183.098862
Rwneg83_45 in83 sn45 11140.846016
Rwneg83_46 in83 sn46 11140.846016
Rwneg83_47 in83 sn47 11140.846016
Rwneg83_48 in83 sn48 11140.846016
Rwneg83_49 in83 sn49 11140.846016
Rwneg83_50 in83 sn50 11140.846016
Rwneg83_51 in83 sn51 11140.846016
Rwneg83_52 in83 sn52 3183.098862
Rwneg83_53 in83 sn53 11140.846016
Rwneg83_54 in83 sn54 3183.098862
Rwneg83_55 in83 sn55 11140.846016
Rwneg83_56 in83 sn56 3183.098862
Rwneg83_57 in83 sn57 11140.846016
Rwneg83_58 in83 sn58 3183.098862
Rwneg83_59 in83 sn59 3183.098862
Rwneg83_60 in83 sn60 3183.098862
Rwneg83_61 in83 sn61 3183.098862
Rwneg83_62 in83 sn62 11140.846016
Rwneg83_63 in83 sn63 3183.098862
Rwneg83_64 in83 sn64 11140.846016
Rwneg83_65 in83 sn65 11140.846016
Rwneg83_66 in83 sn66 3183.098862
Rwneg83_67 in83 sn67 11140.846016
Rwneg83_68 in83 sn68 11140.846016
Rwneg83_69 in83 sn69 11140.846016
Rwneg83_70 in83 sn70 3183.098862
Rwneg83_71 in83 sn71 11140.846016
Rwneg83_72 in83 sn72 3183.098862
Rwneg83_73 in83 sn73 11140.846016
Rwneg83_74 in83 sn74 11140.846016
Rwneg83_75 in83 sn75 11140.846016
Rwneg83_76 in83 sn76 3183.098862
Rwneg83_77 in83 sn77 11140.846016
Rwneg83_78 in83 sn78 11140.846016
Rwneg83_79 in83 sn79 3183.098862
Rwneg83_80 in83 sn80 11140.846016
Rwneg83_81 in83 sn81 11140.846016
Rwneg83_82 in83 sn82 3183.098862
Rwneg83_83 in83 sn83 11140.846016
Rwneg83_84 in83 sn84 3183.098862
Rwneg83_85 in83 sn85 11140.846016
Rwneg83_86 in83 sn86 3183.098862
Rwneg83_87 in83 sn87 11140.846016
Rwneg83_88 in83 sn88 3183.098862
Rwneg83_89 in83 sn89 11140.846016
Rwneg83_90 in83 sn90 11140.846016
Rwneg83_91 in83 sn91 3183.098862
Rwneg83_92 in83 sn92 3183.098862
Rwneg83_93 in83 sn93 11140.846016
Rwneg83_94 in83 sn94 11140.846016
Rwneg83_95 in83 sn95 11140.846016
Rwneg83_96 in83 sn96 3183.098862
Rwneg83_97 in83 sn97 11140.846016
Rwneg83_98 in83 sn98 11140.846016
Rwneg83_99 in83 sn99 11140.846016
Rwneg83_100 in83 sn100 11140.846016
Rwneg84_1 in84 sn1 11140.846016
Rwneg84_2 in84 sn2 3183.098862
Rwneg84_3 in84 sn3 3183.098862
Rwneg84_4 in84 sn4 3183.098862
Rwneg84_5 in84 sn5 11140.846016
Rwneg84_6 in84 sn6 3183.098862
Rwneg84_7 in84 sn7 11140.846016
Rwneg84_8 in84 sn8 11140.846016
Rwneg84_9 in84 sn9 11140.846016
Rwneg84_10 in84 sn10 11140.846016
Rwneg84_11 in84 sn11 11140.846016
Rwneg84_12 in84 sn12 3183.098862
Rwneg84_13 in84 sn13 11140.846016
Rwneg84_14 in84 sn14 11140.846016
Rwneg84_15 in84 sn15 3183.098862
Rwneg84_16 in84 sn16 11140.846016
Rwneg84_17 in84 sn17 11140.846016
Rwneg84_18 in84 sn18 11140.846016
Rwneg84_19 in84 sn19 11140.846016
Rwneg84_20 in84 sn20 3183.098862
Rwneg84_21 in84 sn21 11140.846016
Rwneg84_22 in84 sn22 11140.846016
Rwneg84_23 in84 sn23 11140.846016
Rwneg84_24 in84 sn24 11140.846016
Rwneg84_25 in84 sn25 11140.846016
Rwneg84_26 in84 sn26 3183.098862
Rwneg84_27 in84 sn27 3183.098862
Rwneg84_28 in84 sn28 11140.846016
Rwneg84_29 in84 sn29 3183.098862
Rwneg84_30 in84 sn30 11140.846016
Rwneg84_31 in84 sn31 3183.098862
Rwneg84_32 in84 sn32 3183.098862
Rwneg84_33 in84 sn33 11140.846016
Rwneg84_34 in84 sn34 11140.846016
Rwneg84_35 in84 sn35 11140.846016
Rwneg84_36 in84 sn36 3183.098862
Rwneg84_37 in84 sn37 11140.846016
Rwneg84_38 in84 sn38 11140.846016
Rwneg84_39 in84 sn39 11140.846016
Rwneg84_40 in84 sn40 11140.846016
Rwneg84_41 in84 sn41 11140.846016
Rwneg84_42 in84 sn42 3183.098862
Rwneg84_43 in84 sn43 3183.098862
Rwneg84_44 in84 sn44 11140.846016
Rwneg84_45 in84 sn45 3183.098862
Rwneg84_46 in84 sn46 3183.098862
Rwneg84_47 in84 sn47 3183.098862
Rwneg84_48 in84 sn48 11140.846016
Rwneg84_49 in84 sn49 3183.098862
Rwneg84_50 in84 sn50 11140.846016
Rwneg84_51 in84 sn51 11140.846016
Rwneg84_52 in84 sn52 3183.098862
Rwneg84_53 in84 sn53 3183.098862
Rwneg84_54 in84 sn54 11140.846016
Rwneg84_55 in84 sn55 3183.098862
Rwneg84_56 in84 sn56 11140.846016
Rwneg84_57 in84 sn57 3183.098862
Rwneg84_58 in84 sn58 3183.098862
Rwneg84_59 in84 sn59 3183.098862
Rwneg84_60 in84 sn60 11140.846016
Rwneg84_61 in84 sn61 3183.098862
Rwneg84_62 in84 sn62 11140.846016
Rwneg84_63 in84 sn63 11140.846016
Rwneg84_64 in84 sn64 3183.098862
Rwneg84_65 in84 sn65 11140.846016
Rwneg84_66 in84 sn66 11140.846016
Rwneg84_67 in84 sn67 11140.846016
Rwneg84_68 in84 sn68 3183.098862
Rwneg84_69 in84 sn69 11140.846016
Rwneg84_70 in84 sn70 11140.846016
Rwneg84_71 in84 sn71 11140.846016
Rwneg84_72 in84 sn72 11140.846016
Rwneg84_73 in84 sn73 3183.098862
Rwneg84_74 in84 sn74 3183.098862
Rwneg84_75 in84 sn75 11140.846016
Rwneg84_76 in84 sn76 11140.846016
Rwneg84_77 in84 sn77 11140.846016
Rwneg84_78 in84 sn78 11140.846016
Rwneg84_79 in84 sn79 3183.098862
Rwneg84_80 in84 sn80 3183.098862
Rwneg84_81 in84 sn81 11140.846016
Rwneg84_82 in84 sn82 11140.846016
Rwneg84_83 in84 sn83 11140.846016
Rwneg84_84 in84 sn84 3183.098862
Rwneg84_85 in84 sn85 11140.846016
Rwneg84_86 in84 sn86 11140.846016
Rwneg84_87 in84 sn87 11140.846016
Rwneg84_88 in84 sn88 11140.846016
Rwneg84_89 in84 sn89 11140.846016
Rwneg84_90 in84 sn90 3183.098862
Rwneg84_91 in84 sn91 11140.846016
Rwneg84_92 in84 sn92 11140.846016
Rwneg84_93 in84 sn93 3183.098862
Rwneg84_94 in84 sn94 11140.846016
Rwneg84_95 in84 sn95 11140.846016
Rwneg84_96 in84 sn96 11140.846016
Rwneg84_97 in84 sn97 3183.098862
Rwneg84_98 in84 sn98 11140.846016
Rwneg84_99 in84 sn99 11140.846016
Rwneg84_100 in84 sn100 11140.846016
Rwneg85_1 in85 sn1 3183.098862
Rwneg85_2 in85 sn2 11140.846016
Rwneg85_3 in85 sn3 11140.846016
Rwneg85_4 in85 sn4 11140.846016
Rwneg85_5 in85 sn5 11140.846016
Rwneg85_6 in85 sn6 3183.098862
Rwneg85_7 in85 sn7 11140.846016
Rwneg85_8 in85 sn8 11140.846016
Rwneg85_9 in85 sn9 11140.846016
Rwneg85_10 in85 sn10 11140.846016
Rwneg85_11 in85 sn11 3183.098862
Rwneg85_12 in85 sn12 3183.098862
Rwneg85_13 in85 sn13 11140.846016
Rwneg85_14 in85 sn14 3183.098862
Rwneg85_15 in85 sn15 11140.846016
Rwneg85_16 in85 sn16 3183.098862
Rwneg85_17 in85 sn17 11140.846016
Rwneg85_18 in85 sn18 11140.846016
Rwneg85_19 in85 sn19 3183.098862
Rwneg85_20 in85 sn20 11140.846016
Rwneg85_21 in85 sn21 11140.846016
Rwneg85_22 in85 sn22 3183.098862
Rwneg85_23 in85 sn23 3183.098862
Rwneg85_24 in85 sn24 11140.846016
Rwneg85_25 in85 sn25 3183.098862
Rwneg85_26 in85 sn26 11140.846016
Rwneg85_27 in85 sn27 3183.098862
Rwneg85_28 in85 sn28 3183.098862
Rwneg85_29 in85 sn29 3183.098862
Rwneg85_30 in85 sn30 11140.846016
Rwneg85_31 in85 sn31 11140.846016
Rwneg85_32 in85 sn32 3183.098862
Rwneg85_33 in85 sn33 11140.846016
Rwneg85_34 in85 sn34 11140.846016
Rwneg85_35 in85 sn35 3183.098862
Rwneg85_36 in85 sn36 11140.846016
Rwneg85_37 in85 sn37 11140.846016
Rwneg85_38 in85 sn38 11140.846016
Rwneg85_39 in85 sn39 11140.846016
Rwneg85_40 in85 sn40 11140.846016
Rwneg85_41 in85 sn41 3183.098862
Rwneg85_42 in85 sn42 11140.846016
Rwneg85_43 in85 sn43 3183.098862
Rwneg85_44 in85 sn44 3183.098862
Rwneg85_45 in85 sn45 3183.098862
Rwneg85_46 in85 sn46 11140.846016
Rwneg85_47 in85 sn47 11140.846016
Rwneg85_48 in85 sn48 3183.098862
Rwneg85_49 in85 sn49 11140.846016
Rwneg85_50 in85 sn50 11140.846016
Rwneg85_51 in85 sn51 11140.846016
Rwneg85_52 in85 sn52 11140.846016
Rwneg85_53 in85 sn53 11140.846016
Rwneg85_54 in85 sn54 11140.846016
Rwneg85_55 in85 sn55 3183.098862
Rwneg85_56 in85 sn56 11140.846016
Rwneg85_57 in85 sn57 11140.846016
Rwneg85_58 in85 sn58 11140.846016
Rwneg85_59 in85 sn59 3183.098862
Rwneg85_60 in85 sn60 3183.098862
Rwneg85_61 in85 sn61 3183.098862
Rwneg85_62 in85 sn62 3183.098862
Rwneg85_63 in85 sn63 11140.846016
Rwneg85_64 in85 sn64 3183.098862
Rwneg85_65 in85 sn65 11140.846016
Rwneg85_66 in85 sn66 11140.846016
Rwneg85_67 in85 sn67 11140.846016
Rwneg85_68 in85 sn68 11140.846016
Rwneg85_69 in85 sn69 11140.846016
Rwneg85_70 in85 sn70 11140.846016
Rwneg85_71 in85 sn71 11140.846016
Rwneg85_72 in85 sn72 3183.098862
Rwneg85_73 in85 sn73 3183.098862
Rwneg85_74 in85 sn74 3183.098862
Rwneg85_75 in85 sn75 3183.098862
Rwneg85_76 in85 sn76 3183.098862
Rwneg85_77 in85 sn77 3183.098862
Rwneg85_78 in85 sn78 11140.846016
Rwneg85_79 in85 sn79 11140.846016
Rwneg85_80 in85 sn80 3183.098862
Rwneg85_81 in85 sn81 11140.846016
Rwneg85_82 in85 sn82 11140.846016
Rwneg85_83 in85 sn83 11140.846016
Rwneg85_84 in85 sn84 3183.098862
Rwneg85_85 in85 sn85 11140.846016
Rwneg85_86 in85 sn86 3183.098862
Rwneg85_87 in85 sn87 3183.098862
Rwneg85_88 in85 sn88 11140.846016
Rwneg85_89 in85 sn89 3183.098862
Rwneg85_90 in85 sn90 11140.846016
Rwneg85_91 in85 sn91 3183.098862
Rwneg85_92 in85 sn92 11140.846016
Rwneg85_93 in85 sn93 11140.846016
Rwneg85_94 in85 sn94 3183.098862
Rwneg85_95 in85 sn95 3183.098862
Rwneg85_96 in85 sn96 11140.846016
Rwneg85_97 in85 sn97 11140.846016
Rwneg85_98 in85 sn98 11140.846016
Rwneg85_99 in85 sn99 11140.846016
Rwneg85_100 in85 sn100 11140.846016
Rwneg86_1 in86 sn1 11140.846016
Rwneg86_2 in86 sn2 3183.098862
Rwneg86_3 in86 sn3 11140.846016
Rwneg86_4 in86 sn4 3183.098862
Rwneg86_5 in86 sn5 11140.846016
Rwneg86_6 in86 sn6 11140.846016
Rwneg86_7 in86 sn7 11140.846016
Rwneg86_8 in86 sn8 11140.846016
Rwneg86_9 in86 sn9 3183.098862
Rwneg86_10 in86 sn10 11140.846016
Rwneg86_11 in86 sn11 11140.846016
Rwneg86_12 in86 sn12 3183.098862
Rwneg86_13 in86 sn13 11140.846016
Rwneg86_14 in86 sn14 11140.846016
Rwneg86_15 in86 sn15 3183.098862
Rwneg86_16 in86 sn16 11140.846016
Rwneg86_17 in86 sn17 11140.846016
Rwneg86_18 in86 sn18 3183.098862
Rwneg86_19 in86 sn19 11140.846016
Rwneg86_20 in86 sn20 11140.846016
Rwneg86_21 in86 sn21 3183.098862
Rwneg86_22 in86 sn22 11140.846016
Rwneg86_23 in86 sn23 11140.846016
Rwneg86_24 in86 sn24 3183.098862
Rwneg86_25 in86 sn25 11140.846016
Rwneg86_26 in86 sn26 3183.098862
Rwneg86_27 in86 sn27 11140.846016
Rwneg86_28 in86 sn28 11140.846016
Rwneg86_29 in86 sn29 3183.098862
Rwneg86_30 in86 sn30 11140.846016
Rwneg86_31 in86 sn31 3183.098862
Rwneg86_32 in86 sn32 11140.846016
Rwneg86_33 in86 sn33 11140.846016
Rwneg86_34 in86 sn34 3183.098862
Rwneg86_35 in86 sn35 3183.098862
Rwneg86_36 in86 sn36 3183.098862
Rwneg86_37 in86 sn37 11140.846016
Rwneg86_38 in86 sn38 11140.846016
Rwneg86_39 in86 sn39 3183.098862
Rwneg86_40 in86 sn40 3183.098862
Rwneg86_41 in86 sn41 3183.098862
Rwneg86_42 in86 sn42 3183.098862
Rwneg86_43 in86 sn43 3183.098862
Rwneg86_44 in86 sn44 3183.098862
Rwneg86_45 in86 sn45 3183.098862
Rwneg86_46 in86 sn46 3183.098862
Rwneg86_47 in86 sn47 11140.846016
Rwneg86_48 in86 sn48 3183.098862
Rwneg86_49 in86 sn49 3183.098862
Rwneg86_50 in86 sn50 3183.098862
Rwneg86_51 in86 sn51 3183.098862
Rwneg86_52 in86 sn52 11140.846016
Rwneg86_53 in86 sn53 3183.098862
Rwneg86_54 in86 sn54 3183.098862
Rwneg86_55 in86 sn55 11140.846016
Rwneg86_56 in86 sn56 11140.846016
Rwneg86_57 in86 sn57 11140.846016
Rwneg86_58 in86 sn58 11140.846016
Rwneg86_59 in86 sn59 3183.098862
Rwneg86_60 in86 sn60 3183.098862
Rwneg86_61 in86 sn61 3183.098862
Rwneg86_62 in86 sn62 3183.098862
Rwneg86_63 in86 sn63 3183.098862
Rwneg86_64 in86 sn64 11140.846016
Rwneg86_65 in86 sn65 11140.846016
Rwneg86_66 in86 sn66 3183.098862
Rwneg86_67 in86 sn67 11140.846016
Rwneg86_68 in86 sn68 11140.846016
Rwneg86_69 in86 sn69 3183.098862
Rwneg86_70 in86 sn70 3183.098862
Rwneg86_71 in86 sn71 3183.098862
Rwneg86_72 in86 sn72 3183.098862
Rwneg86_73 in86 sn73 11140.846016
Rwneg86_74 in86 sn74 3183.098862
Rwneg86_75 in86 sn75 11140.846016
Rwneg86_76 in86 sn76 11140.846016
Rwneg86_77 in86 sn77 3183.098862
Rwneg86_78 in86 sn78 11140.846016
Rwneg86_79 in86 sn79 11140.846016
Rwneg86_80 in86 sn80 11140.846016
Rwneg86_81 in86 sn81 3183.098862
Rwneg86_82 in86 sn82 3183.098862
Rwneg86_83 in86 sn83 11140.846016
Rwneg86_84 in86 sn84 11140.846016
Rwneg86_85 in86 sn85 3183.098862
Rwneg86_86 in86 sn86 11140.846016
Rwneg86_87 in86 sn87 3183.098862
Rwneg86_88 in86 sn88 11140.846016
Rwneg86_89 in86 sn89 3183.098862
Rwneg86_90 in86 sn90 11140.846016
Rwneg86_91 in86 sn91 11140.846016
Rwneg86_92 in86 sn92 3183.098862
Rwneg86_93 in86 sn93 3183.098862
Rwneg86_94 in86 sn94 11140.846016
Rwneg86_95 in86 sn95 11140.846016
Rwneg86_96 in86 sn96 11140.846016
Rwneg86_97 in86 sn97 11140.846016
Rwneg86_98 in86 sn98 3183.098862
Rwneg86_99 in86 sn99 3183.098862
Rwneg86_100 in86 sn100 11140.846016
Rwneg87_1 in87 sn1 11140.846016
Rwneg87_2 in87 sn2 11140.846016
Rwneg87_3 in87 sn3 3183.098862
Rwneg87_4 in87 sn4 3183.098862
Rwneg87_5 in87 sn5 3183.098862
Rwneg87_6 in87 sn6 11140.846016
Rwneg87_7 in87 sn7 11140.846016
Rwneg87_8 in87 sn8 3183.098862
Rwneg87_9 in87 sn9 11140.846016
Rwneg87_10 in87 sn10 11140.846016
Rwneg87_11 in87 sn11 11140.846016
Rwneg87_12 in87 sn12 11140.846016
Rwneg87_13 in87 sn13 3183.098862
Rwneg87_14 in87 sn14 11140.846016
Rwneg87_15 in87 sn15 3183.098862
Rwneg87_16 in87 sn16 11140.846016
Rwneg87_17 in87 sn17 3183.098862
Rwneg87_18 in87 sn18 11140.846016
Rwneg87_19 in87 sn19 3183.098862
Rwneg87_20 in87 sn20 3183.098862
Rwneg87_21 in87 sn21 3183.098862
Rwneg87_22 in87 sn22 11140.846016
Rwneg87_23 in87 sn23 11140.846016
Rwneg87_24 in87 sn24 11140.846016
Rwneg87_25 in87 sn25 11140.846016
Rwneg87_26 in87 sn26 11140.846016
Rwneg87_27 in87 sn27 11140.846016
Rwneg87_28 in87 sn28 11140.846016
Rwneg87_29 in87 sn29 3183.098862
Rwneg87_30 in87 sn30 11140.846016
Rwneg87_31 in87 sn31 11140.846016
Rwneg87_32 in87 sn32 11140.846016
Rwneg87_33 in87 sn33 11140.846016
Rwneg87_34 in87 sn34 11140.846016
Rwneg87_35 in87 sn35 11140.846016
Rwneg87_36 in87 sn36 3183.098862
Rwneg87_37 in87 sn37 3183.098862
Rwneg87_38 in87 sn38 3183.098862
Rwneg87_39 in87 sn39 11140.846016
Rwneg87_40 in87 sn40 3183.098862
Rwneg87_41 in87 sn41 11140.846016
Rwneg87_42 in87 sn42 3183.098862
Rwneg87_43 in87 sn43 11140.846016
Rwneg87_44 in87 sn44 11140.846016
Rwneg87_45 in87 sn45 11140.846016
Rwneg87_46 in87 sn46 11140.846016
Rwneg87_47 in87 sn47 3183.098862
Rwneg87_48 in87 sn48 11140.846016
Rwneg87_49 in87 sn49 3183.098862
Rwneg87_50 in87 sn50 11140.846016
Rwneg87_51 in87 sn51 3183.098862
Rwneg87_52 in87 sn52 11140.846016
Rwneg87_53 in87 sn53 3183.098862
Rwneg87_54 in87 sn54 3183.098862
Rwneg87_55 in87 sn55 3183.098862
Rwneg87_56 in87 sn56 3183.098862
Rwneg87_57 in87 sn57 11140.846016
Rwneg87_58 in87 sn58 3183.098862
Rwneg87_59 in87 sn59 11140.846016
Rwneg87_60 in87 sn60 3183.098862
Rwneg87_61 in87 sn61 3183.098862
Rwneg87_62 in87 sn62 11140.846016
Rwneg87_63 in87 sn63 3183.098862
Rwneg87_64 in87 sn64 11140.846016
Rwneg87_65 in87 sn65 3183.098862
Rwneg87_66 in87 sn66 3183.098862
Rwneg87_67 in87 sn67 11140.846016
Rwneg87_68 in87 sn68 3183.098862
Rwneg87_69 in87 sn69 3183.098862
Rwneg87_70 in87 sn70 3183.098862
Rwneg87_71 in87 sn71 3183.098862
Rwneg87_72 in87 sn72 3183.098862
Rwneg87_73 in87 sn73 11140.846016
Rwneg87_74 in87 sn74 3183.098862
Rwneg87_75 in87 sn75 11140.846016
Rwneg87_76 in87 sn76 11140.846016
Rwneg87_77 in87 sn77 3183.098862
Rwneg87_78 in87 sn78 3183.098862
Rwneg87_79 in87 sn79 3183.098862
Rwneg87_80 in87 sn80 11140.846016
Rwneg87_81 in87 sn81 11140.846016
Rwneg87_82 in87 sn82 3183.098862
Rwneg87_83 in87 sn83 11140.846016
Rwneg87_84 in87 sn84 3183.098862
Rwneg87_85 in87 sn85 3183.098862
Rwneg87_86 in87 sn86 3183.098862
Rwneg87_87 in87 sn87 3183.098862
Rwneg87_88 in87 sn88 3183.098862
Rwneg87_89 in87 sn89 11140.846016
Rwneg87_90 in87 sn90 3183.098862
Rwneg87_91 in87 sn91 11140.846016
Rwneg87_92 in87 sn92 11140.846016
Rwneg87_93 in87 sn93 11140.846016
Rwneg87_94 in87 sn94 3183.098862
Rwneg87_95 in87 sn95 11140.846016
Rwneg87_96 in87 sn96 11140.846016
Rwneg87_97 in87 sn97 11140.846016
Rwneg87_98 in87 sn98 3183.098862
Rwneg87_99 in87 sn99 11140.846016
Rwneg87_100 in87 sn100 3183.098862
Rwneg88_1 in88 sn1 11140.846016
Rwneg88_2 in88 sn2 3183.098862
Rwneg88_3 in88 sn3 3183.098862
Rwneg88_4 in88 sn4 3183.098862
Rwneg88_5 in88 sn5 11140.846016
Rwneg88_6 in88 sn6 11140.846016
Rwneg88_7 in88 sn7 11140.846016
Rwneg88_8 in88 sn8 3183.098862
Rwneg88_9 in88 sn9 3183.098862
Rwneg88_10 in88 sn10 3183.098862
Rwneg88_11 in88 sn11 11140.846016
Rwneg88_12 in88 sn12 11140.846016
Rwneg88_13 in88 sn13 11140.846016
Rwneg88_14 in88 sn14 11140.846016
Rwneg88_15 in88 sn15 11140.846016
Rwneg88_16 in88 sn16 3183.098862
Rwneg88_17 in88 sn17 3183.098862
Rwneg88_18 in88 sn18 3183.098862
Rwneg88_19 in88 sn19 11140.846016
Rwneg88_20 in88 sn20 3183.098862
Rwneg88_21 in88 sn21 11140.846016
Rwneg88_22 in88 sn22 11140.846016
Rwneg88_23 in88 sn23 11140.846016
Rwneg88_24 in88 sn24 3183.098862
Rwneg88_25 in88 sn25 3183.098862
Rwneg88_26 in88 sn26 11140.846016
Rwneg88_27 in88 sn27 3183.098862
Rwneg88_28 in88 sn28 11140.846016
Rwneg88_29 in88 sn29 11140.846016
Rwneg88_30 in88 sn30 3183.098862
Rwneg88_31 in88 sn31 3183.098862
Rwneg88_32 in88 sn32 3183.098862
Rwneg88_33 in88 sn33 11140.846016
Rwneg88_34 in88 sn34 11140.846016
Rwneg88_35 in88 sn35 3183.098862
Rwneg88_36 in88 sn36 3183.098862
Rwneg88_37 in88 sn37 11140.846016
Rwneg88_38 in88 sn38 11140.846016
Rwneg88_39 in88 sn39 11140.846016
Rwneg88_40 in88 sn40 11140.846016
Rwneg88_41 in88 sn41 3183.098862
Rwneg88_42 in88 sn42 11140.846016
Rwneg88_43 in88 sn43 3183.098862
Rwneg88_44 in88 sn44 11140.846016
Rwneg88_45 in88 sn45 3183.098862
Rwneg88_46 in88 sn46 11140.846016
Rwneg88_47 in88 sn47 11140.846016
Rwneg88_48 in88 sn48 3183.098862
Rwneg88_49 in88 sn49 11140.846016
Rwneg88_50 in88 sn50 11140.846016
Rwneg88_51 in88 sn51 11140.846016
Rwneg88_52 in88 sn52 3183.098862
Rwneg88_53 in88 sn53 11140.846016
Rwneg88_54 in88 sn54 11140.846016
Rwneg88_55 in88 sn55 11140.846016
Rwneg88_56 in88 sn56 3183.098862
Rwneg88_57 in88 sn57 3183.098862
Rwneg88_58 in88 sn58 11140.846016
Rwneg88_59 in88 sn59 3183.098862
Rwneg88_60 in88 sn60 3183.098862
Rwneg88_61 in88 sn61 11140.846016
Rwneg88_62 in88 sn62 3183.098862
Rwneg88_63 in88 sn63 11140.846016
Rwneg88_64 in88 sn64 11140.846016
Rwneg88_65 in88 sn65 3183.098862
Rwneg88_66 in88 sn66 11140.846016
Rwneg88_67 in88 sn67 11140.846016
Rwneg88_68 in88 sn68 3183.098862
Rwneg88_69 in88 sn69 3183.098862
Rwneg88_70 in88 sn70 11140.846016
Rwneg88_71 in88 sn71 11140.846016
Rwneg88_72 in88 sn72 11140.846016
Rwneg88_73 in88 sn73 3183.098862
Rwneg88_74 in88 sn74 3183.098862
Rwneg88_75 in88 sn75 11140.846016
Rwneg88_76 in88 sn76 11140.846016
Rwneg88_77 in88 sn77 3183.098862
Rwneg88_78 in88 sn78 11140.846016
Rwneg88_79 in88 sn79 3183.098862
Rwneg88_80 in88 sn80 3183.098862
Rwneg88_81 in88 sn81 3183.098862
Rwneg88_82 in88 sn82 11140.846016
Rwneg88_83 in88 sn83 3183.098862
Rwneg88_84 in88 sn84 3183.098862
Rwneg88_85 in88 sn85 3183.098862
Rwneg88_86 in88 sn86 11140.846016
Rwneg88_87 in88 sn87 11140.846016
Rwneg88_88 in88 sn88 11140.846016
Rwneg88_89 in88 sn89 11140.846016
Rwneg88_90 in88 sn90 3183.098862
Rwneg88_91 in88 sn91 3183.098862
Rwneg88_92 in88 sn92 3183.098862
Rwneg88_93 in88 sn93 11140.846016
Rwneg88_94 in88 sn94 3183.098862
Rwneg88_95 in88 sn95 3183.098862
Rwneg88_96 in88 sn96 3183.098862
Rwneg88_97 in88 sn97 11140.846016
Rwneg88_98 in88 sn98 3183.098862
Rwneg88_99 in88 sn99 11140.846016
Rwneg88_100 in88 sn100 11140.846016
Rwneg89_1 in89 sn1 11140.846016
Rwneg89_2 in89 sn2 11140.846016
Rwneg89_3 in89 sn3 11140.846016
Rwneg89_4 in89 sn4 11140.846016
Rwneg89_5 in89 sn5 3183.098862
Rwneg89_6 in89 sn6 3183.098862
Rwneg89_7 in89 sn7 3183.098862
Rwneg89_8 in89 sn8 11140.846016
Rwneg89_9 in89 sn9 11140.846016
Rwneg89_10 in89 sn10 3183.098862
Rwneg89_11 in89 sn11 3183.098862
Rwneg89_12 in89 sn12 11140.846016
Rwneg89_13 in89 sn13 11140.846016
Rwneg89_14 in89 sn14 11140.846016
Rwneg89_15 in89 sn15 11140.846016
Rwneg89_16 in89 sn16 3183.098862
Rwneg89_17 in89 sn17 3183.098862
Rwneg89_18 in89 sn18 11140.846016
Rwneg89_19 in89 sn19 11140.846016
Rwneg89_20 in89 sn20 11140.846016
Rwneg89_21 in89 sn21 3183.098862
Rwneg89_22 in89 sn22 3183.098862
Rwneg89_23 in89 sn23 11140.846016
Rwneg89_24 in89 sn24 11140.846016
Rwneg89_25 in89 sn25 3183.098862
Rwneg89_26 in89 sn26 3183.098862
Rwneg89_27 in89 sn27 3183.098862
Rwneg89_28 in89 sn28 3183.098862
Rwneg89_29 in89 sn29 3183.098862
Rwneg89_30 in89 sn30 11140.846016
Rwneg89_31 in89 sn31 11140.846016
Rwneg89_32 in89 sn32 11140.846016
Rwneg89_33 in89 sn33 3183.098862
Rwneg89_34 in89 sn34 11140.846016
Rwneg89_35 in89 sn35 3183.098862
Rwneg89_36 in89 sn36 11140.846016
Rwneg89_37 in89 sn37 3183.098862
Rwneg89_38 in89 sn38 3183.098862
Rwneg89_39 in89 sn39 3183.098862
Rwneg89_40 in89 sn40 11140.846016
Rwneg89_41 in89 sn41 11140.846016
Rwneg89_42 in89 sn42 11140.846016
Rwneg89_43 in89 sn43 3183.098862
Rwneg89_44 in89 sn44 11140.846016
Rwneg89_45 in89 sn45 11140.846016
Rwneg89_46 in89 sn46 3183.098862
Rwneg89_47 in89 sn47 11140.846016
Rwneg89_48 in89 sn48 3183.098862
Rwneg89_49 in89 sn49 11140.846016
Rwneg89_50 in89 sn50 11140.846016
Rwneg89_51 in89 sn51 11140.846016
Rwneg89_52 in89 sn52 11140.846016
Rwneg89_53 in89 sn53 3183.098862
Rwneg89_54 in89 sn54 3183.098862
Rwneg89_55 in89 sn55 3183.098862
Rwneg89_56 in89 sn56 11140.846016
Rwneg89_57 in89 sn57 11140.846016
Rwneg89_58 in89 sn58 11140.846016
Rwneg89_59 in89 sn59 3183.098862
Rwneg89_60 in89 sn60 3183.098862
Rwneg89_61 in89 sn61 3183.098862
Rwneg89_62 in89 sn62 11140.846016
Rwneg89_63 in89 sn63 11140.846016
Rwneg89_64 in89 sn64 3183.098862
Rwneg89_65 in89 sn65 3183.098862
Rwneg89_66 in89 sn66 11140.846016
Rwneg89_67 in89 sn67 3183.098862
Rwneg89_68 in89 sn68 11140.846016
Rwneg89_69 in89 sn69 11140.846016
Rwneg89_70 in89 sn70 11140.846016
Rwneg89_71 in89 sn71 11140.846016
Rwneg89_72 in89 sn72 11140.846016
Rwneg89_73 in89 sn73 3183.098862
Rwneg89_74 in89 sn74 11140.846016
Rwneg89_75 in89 sn75 3183.098862
Rwneg89_76 in89 sn76 3183.098862
Rwneg89_77 in89 sn77 3183.098862
Rwneg89_78 in89 sn78 11140.846016
Rwneg89_79 in89 sn79 11140.846016
Rwneg89_80 in89 sn80 3183.098862
Rwneg89_81 in89 sn81 3183.098862
Rwneg89_82 in89 sn82 11140.846016
Rwneg89_83 in89 sn83 11140.846016
Rwneg89_84 in89 sn84 11140.846016
Rwneg89_85 in89 sn85 11140.846016
Rwneg89_86 in89 sn86 11140.846016
Rwneg89_87 in89 sn87 11140.846016
Rwneg89_88 in89 sn88 11140.846016
Rwneg89_89 in89 sn89 3183.098862
Rwneg89_90 in89 sn90 11140.846016
Rwneg89_91 in89 sn91 3183.098862
Rwneg89_92 in89 sn92 3183.098862
Rwneg89_93 in89 sn93 11140.846016
Rwneg89_94 in89 sn94 3183.098862
Rwneg89_95 in89 sn95 11140.846016
Rwneg89_96 in89 sn96 3183.098862
Rwneg89_97 in89 sn97 11140.846016
Rwneg89_98 in89 sn98 11140.846016
Rwneg89_99 in89 sn99 11140.846016
Rwneg89_100 in89 sn100 3183.098862
Rwneg90_1 in90 sn1 11140.846016
Rwneg90_2 in90 sn2 11140.846016
Rwneg90_3 in90 sn3 11140.846016
Rwneg90_4 in90 sn4 3183.098862
Rwneg90_5 in90 sn5 3183.098862
Rwneg90_6 in90 sn6 11140.846016
Rwneg90_7 in90 sn7 3183.098862
Rwneg90_8 in90 sn8 3183.098862
Rwneg90_9 in90 sn9 3183.098862
Rwneg90_10 in90 sn10 11140.846016
Rwneg90_11 in90 sn11 3183.098862
Rwneg90_12 in90 sn12 3183.098862
Rwneg90_13 in90 sn13 3183.098862
Rwneg90_14 in90 sn14 11140.846016
Rwneg90_15 in90 sn15 11140.846016
Rwneg90_16 in90 sn16 3183.098862
Rwneg90_17 in90 sn17 3183.098862
Rwneg90_18 in90 sn18 11140.846016
Rwneg90_19 in90 sn19 11140.846016
Rwneg90_20 in90 sn20 11140.846016
Rwneg90_21 in90 sn21 3183.098862
Rwneg90_22 in90 sn22 11140.846016
Rwneg90_23 in90 sn23 3183.098862
Rwneg90_24 in90 sn24 11140.846016
Rwneg90_25 in90 sn25 11140.846016
Rwneg90_26 in90 sn26 11140.846016
Rwneg90_27 in90 sn27 3183.098862
Rwneg90_28 in90 sn28 3183.098862
Rwneg90_29 in90 sn29 3183.098862
Rwneg90_30 in90 sn30 3183.098862
Rwneg90_31 in90 sn31 3183.098862
Rwneg90_32 in90 sn32 3183.098862
Rwneg90_33 in90 sn33 3183.098862
Rwneg90_34 in90 sn34 11140.846016
Rwneg90_35 in90 sn35 11140.846016
Rwneg90_36 in90 sn36 11140.846016
Rwneg90_37 in90 sn37 3183.098862
Rwneg90_38 in90 sn38 3183.098862
Rwneg90_39 in90 sn39 3183.098862
Rwneg90_40 in90 sn40 3183.098862
Rwneg90_41 in90 sn41 3183.098862
Rwneg90_42 in90 sn42 11140.846016
Rwneg90_43 in90 sn43 3183.098862
Rwneg90_44 in90 sn44 3183.098862
Rwneg90_45 in90 sn45 3183.098862
Rwneg90_46 in90 sn46 3183.098862
Rwneg90_47 in90 sn47 3183.098862
Rwneg90_48 in90 sn48 11140.846016
Rwneg90_49 in90 sn49 11140.846016
Rwneg90_50 in90 sn50 11140.846016
Rwneg90_51 in90 sn51 3183.098862
Rwneg90_52 in90 sn52 11140.846016
Rwneg90_53 in90 sn53 3183.098862
Rwneg90_54 in90 sn54 3183.098862
Rwneg90_55 in90 sn55 11140.846016
Rwneg90_56 in90 sn56 3183.098862
Rwneg90_57 in90 sn57 3183.098862
Rwneg90_58 in90 sn58 3183.098862
Rwneg90_59 in90 sn59 3183.098862
Rwneg90_60 in90 sn60 3183.098862
Rwneg90_61 in90 sn61 3183.098862
Rwneg90_62 in90 sn62 11140.846016
Rwneg90_63 in90 sn63 3183.098862
Rwneg90_64 in90 sn64 11140.846016
Rwneg90_65 in90 sn65 3183.098862
Rwneg90_66 in90 sn66 3183.098862
Rwneg90_67 in90 sn67 11140.846016
Rwneg90_68 in90 sn68 11140.846016
Rwneg90_69 in90 sn69 3183.098862
Rwneg90_70 in90 sn70 3183.098862
Rwneg90_71 in90 sn71 3183.098862
Rwneg90_72 in90 sn72 3183.098862
Rwneg90_73 in90 sn73 3183.098862
Rwneg90_74 in90 sn74 3183.098862
Rwneg90_75 in90 sn75 11140.846016
Rwneg90_76 in90 sn76 3183.098862
Rwneg90_77 in90 sn77 11140.846016
Rwneg90_78 in90 sn78 3183.098862
Rwneg90_79 in90 sn79 3183.098862
Rwneg90_80 in90 sn80 3183.098862
Rwneg90_81 in90 sn81 11140.846016
Rwneg90_82 in90 sn82 3183.098862
Rwneg90_83 in90 sn83 3183.098862
Rwneg90_84 in90 sn84 3183.098862
Rwneg90_85 in90 sn85 11140.846016
Rwneg90_86 in90 sn86 3183.098862
Rwneg90_87 in90 sn87 11140.846016
Rwneg90_88 in90 sn88 3183.098862
Rwneg90_89 in90 sn89 3183.098862
Rwneg90_90 in90 sn90 3183.098862
Rwneg90_91 in90 sn91 3183.098862
Rwneg90_92 in90 sn92 11140.846016
Rwneg90_93 in90 sn93 3183.098862
Rwneg90_94 in90 sn94 11140.846016
Rwneg90_95 in90 sn95 11140.846016
Rwneg90_96 in90 sn96 3183.098862
Rwneg90_97 in90 sn97 11140.846016
Rwneg90_98 in90 sn98 11140.846016
Rwneg90_99 in90 sn99 3183.098862
Rwneg90_100 in90 sn100 11140.846016
Rwneg91_1 in91 sn1 3183.098862
Rwneg91_2 in91 sn2 3183.098862
Rwneg91_3 in91 sn3 3183.098862
Rwneg91_4 in91 sn4 11140.846016
Rwneg91_5 in91 sn5 3183.098862
Rwneg91_6 in91 sn6 11140.846016
Rwneg91_7 in91 sn7 3183.098862
Rwneg91_8 in91 sn8 11140.846016
Rwneg91_9 in91 sn9 3183.098862
Rwneg91_10 in91 sn10 3183.098862
Rwneg91_11 in91 sn11 3183.098862
Rwneg91_12 in91 sn12 3183.098862
Rwneg91_13 in91 sn13 3183.098862
Rwneg91_14 in91 sn14 3183.098862
Rwneg91_15 in91 sn15 11140.846016
Rwneg91_16 in91 sn16 11140.846016
Rwneg91_17 in91 sn17 3183.098862
Rwneg91_18 in91 sn18 3183.098862
Rwneg91_19 in91 sn19 3183.098862
Rwneg91_20 in91 sn20 11140.846016
Rwneg91_21 in91 sn21 11140.846016
Rwneg91_22 in91 sn22 11140.846016
Rwneg91_23 in91 sn23 11140.846016
Rwneg91_24 in91 sn24 3183.098862
Rwneg91_25 in91 sn25 3183.098862
Rwneg91_26 in91 sn26 11140.846016
Rwneg91_27 in91 sn27 3183.098862
Rwneg91_28 in91 sn28 11140.846016
Rwneg91_29 in91 sn29 11140.846016
Rwneg91_30 in91 sn30 3183.098862
Rwneg91_31 in91 sn31 3183.098862
Rwneg91_32 in91 sn32 11140.846016
Rwneg91_33 in91 sn33 11140.846016
Rwneg91_34 in91 sn34 11140.846016
Rwneg91_35 in91 sn35 3183.098862
Rwneg91_36 in91 sn36 11140.846016
Rwneg91_37 in91 sn37 11140.846016
Rwneg91_38 in91 sn38 3183.098862
Rwneg91_39 in91 sn39 3183.098862
Rwneg91_40 in91 sn40 3183.098862
Rwneg91_41 in91 sn41 3183.098862
Rwneg91_42 in91 sn42 11140.846016
Rwneg91_43 in91 sn43 11140.846016
Rwneg91_44 in91 sn44 11140.846016
Rwneg91_45 in91 sn45 3183.098862
Rwneg91_46 in91 sn46 11140.846016
Rwneg91_47 in91 sn47 11140.846016
Rwneg91_48 in91 sn48 3183.098862
Rwneg91_49 in91 sn49 11140.846016
Rwneg91_50 in91 sn50 11140.846016
Rwneg91_51 in91 sn51 3183.098862
Rwneg91_52 in91 sn52 3183.098862
Rwneg91_53 in91 sn53 3183.098862
Rwneg91_54 in91 sn54 11140.846016
Rwneg91_55 in91 sn55 11140.846016
Rwneg91_56 in91 sn56 11140.846016
Rwneg91_57 in91 sn57 11140.846016
Rwneg91_58 in91 sn58 11140.846016
Rwneg91_59 in91 sn59 11140.846016
Rwneg91_60 in91 sn60 11140.846016
Rwneg91_61 in91 sn61 3183.098862
Rwneg91_62 in91 sn62 11140.846016
Rwneg91_63 in91 sn63 3183.098862
Rwneg91_64 in91 sn64 11140.846016
Rwneg91_65 in91 sn65 3183.098862
Rwneg91_66 in91 sn66 11140.846016
Rwneg91_67 in91 sn67 3183.098862
Rwneg91_68 in91 sn68 3183.098862
Rwneg91_69 in91 sn69 3183.098862
Rwneg91_70 in91 sn70 11140.846016
Rwneg91_71 in91 sn71 3183.098862
Rwneg91_72 in91 sn72 3183.098862
Rwneg91_73 in91 sn73 3183.098862
Rwneg91_74 in91 sn74 3183.098862
Rwneg91_75 in91 sn75 11140.846016
Rwneg91_76 in91 sn76 11140.846016
Rwneg91_77 in91 sn77 11140.846016
Rwneg91_78 in91 sn78 11140.846016
Rwneg91_79 in91 sn79 3183.098862
Rwneg91_80 in91 sn80 11140.846016
Rwneg91_81 in91 sn81 3183.098862
Rwneg91_82 in91 sn82 11140.846016
Rwneg91_83 in91 sn83 3183.098862
Rwneg91_84 in91 sn84 11140.846016
Rwneg91_85 in91 sn85 3183.098862
Rwneg91_86 in91 sn86 11140.846016
Rwneg91_87 in91 sn87 11140.846016
Rwneg91_88 in91 sn88 3183.098862
Rwneg91_89 in91 sn89 11140.846016
Rwneg91_90 in91 sn90 3183.098862
Rwneg91_91 in91 sn91 11140.846016
Rwneg91_92 in91 sn92 11140.846016
Rwneg91_93 in91 sn93 3183.098862
Rwneg91_94 in91 sn94 11140.846016
Rwneg91_95 in91 sn95 3183.098862
Rwneg91_96 in91 sn96 11140.846016
Rwneg91_97 in91 sn97 3183.098862
Rwneg91_98 in91 sn98 11140.846016
Rwneg91_99 in91 sn99 3183.098862
Rwneg91_100 in91 sn100 3183.098862
Rwneg92_1 in92 sn1 3183.098862
Rwneg92_2 in92 sn2 3183.098862
Rwneg92_3 in92 sn3 11140.846016
Rwneg92_4 in92 sn4 3183.098862
Rwneg92_5 in92 sn5 11140.846016
Rwneg92_6 in92 sn6 11140.846016
Rwneg92_7 in92 sn7 11140.846016
Rwneg92_8 in92 sn8 11140.846016
Rwneg92_9 in92 sn9 3183.098862
Rwneg92_10 in92 sn10 3183.098862
Rwneg92_11 in92 sn11 11140.846016
Rwneg92_12 in92 sn12 11140.846016
Rwneg92_13 in92 sn13 3183.098862
Rwneg92_14 in92 sn14 11140.846016
Rwneg92_15 in92 sn15 11140.846016
Rwneg92_16 in92 sn16 3183.098862
Rwneg92_17 in92 sn17 11140.846016
Rwneg92_18 in92 sn18 3183.098862
Rwneg92_19 in92 sn19 11140.846016
Rwneg92_20 in92 sn20 3183.098862
Rwneg92_21 in92 sn21 11140.846016
Rwneg92_22 in92 sn22 11140.846016
Rwneg92_23 in92 sn23 11140.846016
Rwneg92_24 in92 sn24 3183.098862
Rwneg92_25 in92 sn25 11140.846016
Rwneg92_26 in92 sn26 11140.846016
Rwneg92_27 in92 sn27 11140.846016
Rwneg92_28 in92 sn28 11140.846016
Rwneg92_29 in92 sn29 3183.098862
Rwneg92_30 in92 sn30 11140.846016
Rwneg92_31 in92 sn31 3183.098862
Rwneg92_32 in92 sn32 3183.098862
Rwneg92_33 in92 sn33 3183.098862
Rwneg92_34 in92 sn34 3183.098862
Rwneg92_35 in92 sn35 11140.846016
Rwneg92_36 in92 sn36 3183.098862
Rwneg92_37 in92 sn37 11140.846016
Rwneg92_38 in92 sn38 11140.846016
Rwneg92_39 in92 sn39 11140.846016
Rwneg92_40 in92 sn40 3183.098862
Rwneg92_41 in92 sn41 11140.846016
Rwneg92_42 in92 sn42 3183.098862
Rwneg92_43 in92 sn43 3183.098862
Rwneg92_44 in92 sn44 11140.846016
Rwneg92_45 in92 sn45 3183.098862
Rwneg92_46 in92 sn46 3183.098862
Rwneg92_47 in92 sn47 11140.846016
Rwneg92_48 in92 sn48 3183.098862
Rwneg92_49 in92 sn49 3183.098862
Rwneg92_50 in92 sn50 11140.846016
Rwneg92_51 in92 sn51 3183.098862
Rwneg92_52 in92 sn52 3183.098862
Rwneg92_53 in92 sn53 3183.098862
Rwneg92_54 in92 sn54 11140.846016
Rwneg92_55 in92 sn55 11140.846016
Rwneg92_56 in92 sn56 3183.098862
Rwneg92_57 in92 sn57 11140.846016
Rwneg92_58 in92 sn58 3183.098862
Rwneg92_59 in92 sn59 3183.098862
Rwneg92_60 in92 sn60 11140.846016
Rwneg92_61 in92 sn61 3183.098862
Rwneg92_62 in92 sn62 3183.098862
Rwneg92_63 in92 sn63 11140.846016
Rwneg92_64 in92 sn64 3183.098862
Rwneg92_65 in92 sn65 3183.098862
Rwneg92_66 in92 sn66 3183.098862
Rwneg92_67 in92 sn67 3183.098862
Rwneg92_68 in92 sn68 3183.098862
Rwneg92_69 in92 sn69 11140.846016
Rwneg92_70 in92 sn70 11140.846016
Rwneg92_71 in92 sn71 11140.846016
Rwneg92_72 in92 sn72 3183.098862
Rwneg92_73 in92 sn73 3183.098862
Rwneg92_74 in92 sn74 3183.098862
Rwneg92_75 in92 sn75 11140.846016
Rwneg92_76 in92 sn76 11140.846016
Rwneg92_77 in92 sn77 3183.098862
Rwneg92_78 in92 sn78 3183.098862
Rwneg92_79 in92 sn79 11140.846016
Rwneg92_80 in92 sn80 11140.846016
Rwneg92_81 in92 sn81 11140.846016
Rwneg92_82 in92 sn82 11140.846016
Rwneg92_83 in92 sn83 3183.098862
Rwneg92_84 in92 sn84 11140.846016
Rwneg92_85 in92 sn85 11140.846016
Rwneg92_86 in92 sn86 11140.846016
Rwneg92_87 in92 sn87 11140.846016
Rwneg92_88 in92 sn88 3183.098862
Rwneg92_89 in92 sn89 3183.098862
Rwneg92_90 in92 sn90 3183.098862
Rwneg92_91 in92 sn91 3183.098862
Rwneg92_92 in92 sn92 11140.846016
Rwneg92_93 in92 sn93 11140.846016
Rwneg92_94 in92 sn94 3183.098862
Rwneg92_95 in92 sn95 11140.846016
Rwneg92_96 in92 sn96 11140.846016
Rwneg92_97 in92 sn97 3183.098862
Rwneg92_98 in92 sn98 11140.846016
Rwneg92_99 in92 sn99 3183.098862
Rwneg92_100 in92 sn100 3183.098862
Rwneg93_1 in93 sn1 11140.846016
Rwneg93_2 in93 sn2 11140.846016
Rwneg93_3 in93 sn3 11140.846016
Rwneg93_4 in93 sn4 11140.846016
Rwneg93_5 in93 sn5 11140.846016
Rwneg93_6 in93 sn6 3183.098862
Rwneg93_7 in93 sn7 11140.846016
Rwneg93_8 in93 sn8 11140.846016
Rwneg93_9 in93 sn9 3183.098862
Rwneg93_10 in93 sn10 3183.098862
Rwneg93_11 in93 sn11 3183.098862
Rwneg93_12 in93 sn12 11140.846016
Rwneg93_13 in93 sn13 11140.846016
Rwneg93_14 in93 sn14 11140.846016
Rwneg93_15 in93 sn15 11140.846016
Rwneg93_16 in93 sn16 3183.098862
Rwneg93_17 in93 sn17 11140.846016
Rwneg93_18 in93 sn18 11140.846016
Rwneg93_19 in93 sn19 11140.846016
Rwneg93_20 in93 sn20 11140.846016
Rwneg93_21 in93 sn21 11140.846016
Rwneg93_22 in93 sn22 11140.846016
Rwneg93_23 in93 sn23 11140.846016
Rwneg93_24 in93 sn24 11140.846016
Rwneg93_25 in93 sn25 11140.846016
Rwneg93_26 in93 sn26 3183.098862
Rwneg93_27 in93 sn27 3183.098862
Rwneg93_28 in93 sn28 11140.846016
Rwneg93_29 in93 sn29 11140.846016
Rwneg93_30 in93 sn30 3183.098862
Rwneg93_31 in93 sn31 11140.846016
Rwneg93_32 in93 sn32 3183.098862
Rwneg93_33 in93 sn33 3183.098862
Rwneg93_34 in93 sn34 11140.846016
Rwneg93_35 in93 sn35 11140.846016
Rwneg93_36 in93 sn36 11140.846016
Rwneg93_37 in93 sn37 11140.846016
Rwneg93_38 in93 sn38 3183.098862
Rwneg93_39 in93 sn39 3183.098862
Rwneg93_40 in93 sn40 11140.846016
Rwneg93_41 in93 sn41 3183.098862
Rwneg93_42 in93 sn42 3183.098862
Rwneg93_43 in93 sn43 11140.846016
Rwneg93_44 in93 sn44 3183.098862
Rwneg93_45 in93 sn45 11140.846016
Rwneg93_46 in93 sn46 11140.846016
Rwneg93_47 in93 sn47 11140.846016
Rwneg93_48 in93 sn48 3183.098862
Rwneg93_49 in93 sn49 11140.846016
Rwneg93_50 in93 sn50 11140.846016
Rwneg93_51 in93 sn51 11140.846016
Rwneg93_52 in93 sn52 11140.846016
Rwneg93_53 in93 sn53 11140.846016
Rwneg93_54 in93 sn54 3183.098862
Rwneg93_55 in93 sn55 3183.098862
Rwneg93_56 in93 sn56 11140.846016
Rwneg93_57 in93 sn57 11140.846016
Rwneg93_58 in93 sn58 11140.846016
Rwneg93_59 in93 sn59 3183.098862
Rwneg93_60 in93 sn60 11140.846016
Rwneg93_61 in93 sn61 3183.098862
Rwneg93_62 in93 sn62 3183.098862
Rwneg93_63 in93 sn63 11140.846016
Rwneg93_64 in93 sn64 3183.098862
Rwneg93_65 in93 sn65 11140.846016
Rwneg93_66 in93 sn66 11140.846016
Rwneg93_67 in93 sn67 11140.846016
Rwneg93_68 in93 sn68 11140.846016
Rwneg93_69 in93 sn69 11140.846016
Rwneg93_70 in93 sn70 11140.846016
Rwneg93_71 in93 sn71 3183.098862
Rwneg93_72 in93 sn72 11140.846016
Rwneg93_73 in93 sn73 11140.846016
Rwneg93_74 in93 sn74 11140.846016
Rwneg93_75 in93 sn75 3183.098862
Rwneg93_76 in93 sn76 11140.846016
Rwneg93_77 in93 sn77 11140.846016
Rwneg93_78 in93 sn78 11140.846016
Rwneg93_79 in93 sn79 11140.846016
Rwneg93_80 in93 sn80 3183.098862
Rwneg93_81 in93 sn81 11140.846016
Rwneg93_82 in93 sn82 11140.846016
Rwneg93_83 in93 sn83 11140.846016
Rwneg93_84 in93 sn84 11140.846016
Rwneg93_85 in93 sn85 11140.846016
Rwneg93_86 in93 sn86 3183.098862
Rwneg93_87 in93 sn87 11140.846016
Rwneg93_88 in93 sn88 11140.846016
Rwneg93_89 in93 sn89 3183.098862
Rwneg93_90 in93 sn90 3183.098862
Rwneg93_91 in93 sn91 3183.098862
Rwneg93_92 in93 sn92 3183.098862
Rwneg93_93 in93 sn93 3183.098862
Rwneg93_94 in93 sn94 3183.098862
Rwneg93_95 in93 sn95 11140.846016
Rwneg93_96 in93 sn96 3183.098862
Rwneg93_97 in93 sn97 3183.098862
Rwneg93_98 in93 sn98 11140.846016
Rwneg93_99 in93 sn99 11140.846016
Rwneg93_100 in93 sn100 11140.846016
Rwneg94_1 in94 sn1 11140.846016
Rwneg94_2 in94 sn2 3183.098862
Rwneg94_3 in94 sn3 11140.846016
Rwneg94_4 in94 sn4 11140.846016
Rwneg94_5 in94 sn5 11140.846016
Rwneg94_6 in94 sn6 11140.846016
Rwneg94_7 in94 sn7 11140.846016
Rwneg94_8 in94 sn8 3183.098862
Rwneg94_9 in94 sn9 3183.098862
Rwneg94_10 in94 sn10 3183.098862
Rwneg94_11 in94 sn11 11140.846016
Rwneg94_12 in94 sn12 11140.846016
Rwneg94_13 in94 sn13 11140.846016
Rwneg94_14 in94 sn14 3183.098862
Rwneg94_15 in94 sn15 3183.098862
Rwneg94_16 in94 sn16 11140.846016
Rwneg94_17 in94 sn17 11140.846016
Rwneg94_18 in94 sn18 11140.846016
Rwneg94_19 in94 sn19 11140.846016
Rwneg94_20 in94 sn20 11140.846016
Rwneg94_21 in94 sn21 3183.098862
Rwneg94_22 in94 sn22 11140.846016
Rwneg94_23 in94 sn23 3183.098862
Rwneg94_24 in94 sn24 11140.846016
Rwneg94_25 in94 sn25 3183.098862
Rwneg94_26 in94 sn26 3183.098862
Rwneg94_27 in94 sn27 11140.846016
Rwneg94_28 in94 sn28 3183.098862
Rwneg94_29 in94 sn29 3183.098862
Rwneg94_30 in94 sn30 11140.846016
Rwneg94_31 in94 sn31 11140.846016
Rwneg94_32 in94 sn32 11140.846016
Rwneg94_33 in94 sn33 3183.098862
Rwneg94_34 in94 sn34 11140.846016
Rwneg94_35 in94 sn35 11140.846016
Rwneg94_36 in94 sn36 11140.846016
Rwneg94_37 in94 sn37 11140.846016
Rwneg94_38 in94 sn38 11140.846016
Rwneg94_39 in94 sn39 3183.098862
Rwneg94_40 in94 sn40 3183.098862
Rwneg94_41 in94 sn41 11140.846016
Rwneg94_42 in94 sn42 3183.098862
Rwneg94_43 in94 sn43 11140.846016
Rwneg94_44 in94 sn44 3183.098862
Rwneg94_45 in94 sn45 11140.846016
Rwneg94_46 in94 sn46 11140.846016
Rwneg94_47 in94 sn47 11140.846016
Rwneg94_48 in94 sn48 3183.098862
Rwneg94_49 in94 sn49 3183.098862
Rwneg94_50 in94 sn50 11140.846016
Rwneg94_51 in94 sn51 3183.098862
Rwneg94_52 in94 sn52 3183.098862
Rwneg94_53 in94 sn53 11140.846016
Rwneg94_54 in94 sn54 11140.846016
Rwneg94_55 in94 sn55 3183.098862
Rwneg94_56 in94 sn56 3183.098862
Rwneg94_57 in94 sn57 11140.846016
Rwneg94_58 in94 sn58 3183.098862
Rwneg94_59 in94 sn59 11140.846016
Rwneg94_60 in94 sn60 11140.846016
Rwneg94_61 in94 sn61 11140.846016
Rwneg94_62 in94 sn62 11140.846016
Rwneg94_63 in94 sn63 3183.098862
Rwneg94_64 in94 sn64 3183.098862
Rwneg94_65 in94 sn65 3183.098862
Rwneg94_66 in94 sn66 3183.098862
Rwneg94_67 in94 sn67 3183.098862
Rwneg94_68 in94 sn68 11140.846016
Rwneg94_69 in94 sn69 3183.098862
Rwneg94_70 in94 sn70 3183.098862
Rwneg94_71 in94 sn71 11140.846016
Rwneg94_72 in94 sn72 3183.098862
Rwneg94_73 in94 sn73 11140.846016
Rwneg94_74 in94 sn74 3183.098862
Rwneg94_75 in94 sn75 3183.098862
Rwneg94_76 in94 sn76 11140.846016
Rwneg94_77 in94 sn77 11140.846016
Rwneg94_78 in94 sn78 11140.846016
Rwneg94_79 in94 sn79 3183.098862
Rwneg94_80 in94 sn80 3183.098862
Rwneg94_81 in94 sn81 3183.098862
Rwneg94_82 in94 sn82 3183.098862
Rwneg94_83 in94 sn83 11140.846016
Rwneg94_84 in94 sn84 3183.098862
Rwneg94_85 in94 sn85 11140.846016
Rwneg94_86 in94 sn86 11140.846016
Rwneg94_87 in94 sn87 3183.098862
Rwneg94_88 in94 sn88 3183.098862
Rwneg94_89 in94 sn89 3183.098862
Rwneg94_90 in94 sn90 11140.846016
Rwneg94_91 in94 sn91 3183.098862
Rwneg94_92 in94 sn92 11140.846016
Rwneg94_93 in94 sn93 11140.846016
Rwneg94_94 in94 sn94 11140.846016
Rwneg94_95 in94 sn95 11140.846016
Rwneg94_96 in94 sn96 11140.846016
Rwneg94_97 in94 sn97 11140.846016
Rwneg94_98 in94 sn98 11140.846016
Rwneg94_99 in94 sn99 11140.846016
Rwneg94_100 in94 sn100 11140.846016
Rwneg95_1 in95 sn1 3183.098862
Rwneg95_2 in95 sn2 11140.846016
Rwneg95_3 in95 sn3 3183.098862
Rwneg95_4 in95 sn4 3183.098862
Rwneg95_5 in95 sn5 3183.098862
Rwneg95_6 in95 sn6 11140.846016
Rwneg95_7 in95 sn7 3183.098862
Rwneg95_8 in95 sn8 11140.846016
Rwneg95_9 in95 sn9 11140.846016
Rwneg95_10 in95 sn10 11140.846016
Rwneg95_11 in95 sn11 11140.846016
Rwneg95_12 in95 sn12 3183.098862
Rwneg95_13 in95 sn13 3183.098862
Rwneg95_14 in95 sn14 11140.846016
Rwneg95_15 in95 sn15 11140.846016
Rwneg95_16 in95 sn16 3183.098862
Rwneg95_17 in95 sn17 11140.846016
Rwneg95_18 in95 sn18 11140.846016
Rwneg95_19 in95 sn19 3183.098862
Rwneg95_20 in95 sn20 11140.846016
Rwneg95_21 in95 sn21 11140.846016
Rwneg95_22 in95 sn22 11140.846016
Rwneg95_23 in95 sn23 11140.846016
Rwneg95_24 in95 sn24 11140.846016
Rwneg95_25 in95 sn25 3183.098862
Rwneg95_26 in95 sn26 11140.846016
Rwneg95_27 in95 sn27 11140.846016
Rwneg95_28 in95 sn28 11140.846016
Rwneg95_29 in95 sn29 11140.846016
Rwneg95_30 in95 sn30 3183.098862
Rwneg95_31 in95 sn31 11140.846016
Rwneg95_32 in95 sn32 11140.846016
Rwneg95_33 in95 sn33 3183.098862
Rwneg95_34 in95 sn34 11140.846016
Rwneg95_35 in95 sn35 11140.846016
Rwneg95_36 in95 sn36 3183.098862
Rwneg95_37 in95 sn37 11140.846016
Rwneg95_38 in95 sn38 11140.846016
Rwneg95_39 in95 sn39 11140.846016
Rwneg95_40 in95 sn40 11140.846016
Rwneg95_41 in95 sn41 3183.098862
Rwneg95_42 in95 sn42 11140.846016
Rwneg95_43 in95 sn43 11140.846016
Rwneg95_44 in95 sn44 3183.098862
Rwneg95_45 in95 sn45 11140.846016
Rwneg95_46 in95 sn46 3183.098862
Rwneg95_47 in95 sn47 11140.846016
Rwneg95_48 in95 sn48 3183.098862
Rwneg95_49 in95 sn49 3183.098862
Rwneg95_50 in95 sn50 3183.098862
Rwneg95_51 in95 sn51 3183.098862
Rwneg95_52 in95 sn52 3183.098862
Rwneg95_53 in95 sn53 11140.846016
Rwneg95_54 in95 sn54 11140.846016
Rwneg95_55 in95 sn55 11140.846016
Rwneg95_56 in95 sn56 3183.098862
Rwneg95_57 in95 sn57 3183.098862
Rwneg95_58 in95 sn58 3183.098862
Rwneg95_59 in95 sn59 11140.846016
Rwneg95_60 in95 sn60 3183.098862
Rwneg95_61 in95 sn61 11140.846016
Rwneg95_62 in95 sn62 3183.098862
Rwneg95_63 in95 sn63 11140.846016
Rwneg95_64 in95 sn64 3183.098862
Rwneg95_65 in95 sn65 3183.098862
Rwneg95_66 in95 sn66 11140.846016
Rwneg95_67 in95 sn67 3183.098862
Rwneg95_68 in95 sn68 11140.846016
Rwneg95_69 in95 sn69 11140.846016
Rwneg95_70 in95 sn70 11140.846016
Rwneg95_71 in95 sn71 11140.846016
Rwneg95_72 in95 sn72 11140.846016
Rwneg95_73 in95 sn73 11140.846016
Rwneg95_74 in95 sn74 11140.846016
Rwneg95_75 in95 sn75 11140.846016
Rwneg95_76 in95 sn76 11140.846016
Rwneg95_77 in95 sn77 3183.098862
Rwneg95_78 in95 sn78 3183.098862
Rwneg95_79 in95 sn79 3183.098862
Rwneg95_80 in95 sn80 11140.846016
Rwneg95_81 in95 sn81 11140.846016
Rwneg95_82 in95 sn82 11140.846016
Rwneg95_83 in95 sn83 3183.098862
Rwneg95_84 in95 sn84 3183.098862
Rwneg95_85 in95 sn85 11140.846016
Rwneg95_86 in95 sn86 11140.846016
Rwneg95_87 in95 sn87 11140.846016
Rwneg95_88 in95 sn88 11140.846016
Rwneg95_89 in95 sn89 3183.098862
Rwneg95_90 in95 sn90 11140.846016
Rwneg95_91 in95 sn91 3183.098862
Rwneg95_92 in95 sn92 11140.846016
Rwneg95_93 in95 sn93 3183.098862
Rwneg95_94 in95 sn94 3183.098862
Rwneg95_95 in95 sn95 11140.846016
Rwneg95_96 in95 sn96 11140.846016
Rwneg95_97 in95 sn97 3183.098862
Rwneg95_98 in95 sn98 11140.846016
Rwneg95_99 in95 sn99 3183.098862
Rwneg95_100 in95 sn100 11140.846016
Rwneg96_1 in96 sn1 11140.846016
Rwneg96_2 in96 sn2 3183.098862
Rwneg96_3 in96 sn3 3183.098862
Rwneg96_4 in96 sn4 3183.098862
Rwneg96_5 in96 sn5 3183.098862
Rwneg96_6 in96 sn6 11140.846016
Rwneg96_7 in96 sn7 11140.846016
Rwneg96_8 in96 sn8 11140.846016
Rwneg96_9 in96 sn9 3183.098862
Rwneg96_10 in96 sn10 3183.098862
Rwneg96_11 in96 sn11 11140.846016
Rwneg96_12 in96 sn12 11140.846016
Rwneg96_13 in96 sn13 3183.098862
Rwneg96_14 in96 sn14 11140.846016
Rwneg96_15 in96 sn15 3183.098862
Rwneg96_16 in96 sn16 11140.846016
Rwneg96_17 in96 sn17 3183.098862
Rwneg96_18 in96 sn18 3183.098862
Rwneg96_19 in96 sn19 11140.846016
Rwneg96_20 in96 sn20 11140.846016
Rwneg96_21 in96 sn21 11140.846016
Rwneg96_22 in96 sn22 11140.846016
Rwneg96_23 in96 sn23 11140.846016
Rwneg96_24 in96 sn24 11140.846016
Rwneg96_25 in96 sn25 3183.098862
Rwneg96_26 in96 sn26 3183.098862
Rwneg96_27 in96 sn27 3183.098862
Rwneg96_28 in96 sn28 11140.846016
Rwneg96_29 in96 sn29 3183.098862
Rwneg96_30 in96 sn30 11140.846016
Rwneg96_31 in96 sn31 3183.098862
Rwneg96_32 in96 sn32 3183.098862
Rwneg96_33 in96 sn33 11140.846016
Rwneg96_34 in96 sn34 3183.098862
Rwneg96_35 in96 sn35 11140.846016
Rwneg96_36 in96 sn36 11140.846016
Rwneg96_37 in96 sn37 11140.846016
Rwneg96_38 in96 sn38 11140.846016
Rwneg96_39 in96 sn39 11140.846016
Rwneg96_40 in96 sn40 3183.098862
Rwneg96_41 in96 sn41 11140.846016
Rwneg96_42 in96 sn42 11140.846016
Rwneg96_43 in96 sn43 3183.098862
Rwneg96_44 in96 sn44 11140.846016
Rwneg96_45 in96 sn45 11140.846016
Rwneg96_46 in96 sn46 11140.846016
Rwneg96_47 in96 sn47 3183.098862
Rwneg96_48 in96 sn48 11140.846016
Rwneg96_49 in96 sn49 3183.098862
Rwneg96_50 in96 sn50 3183.098862
Rwneg96_51 in96 sn51 11140.846016
Rwneg96_52 in96 sn52 3183.098862
Rwneg96_53 in96 sn53 11140.846016
Rwneg96_54 in96 sn54 11140.846016
Rwneg96_55 in96 sn55 11140.846016
Rwneg96_56 in96 sn56 11140.846016
Rwneg96_57 in96 sn57 11140.846016
Rwneg96_58 in96 sn58 11140.846016
Rwneg96_59 in96 sn59 3183.098862
Rwneg96_60 in96 sn60 11140.846016
Rwneg96_61 in96 sn61 3183.098862
Rwneg96_62 in96 sn62 11140.846016
Rwneg96_63 in96 sn63 3183.098862
Rwneg96_64 in96 sn64 3183.098862
Rwneg96_65 in96 sn65 3183.098862
Rwneg96_66 in96 sn66 11140.846016
Rwneg96_67 in96 sn67 11140.846016
Rwneg96_68 in96 sn68 3183.098862
Rwneg96_69 in96 sn69 3183.098862
Rwneg96_70 in96 sn70 11140.846016
Rwneg96_71 in96 sn71 11140.846016
Rwneg96_72 in96 sn72 11140.846016
Rwneg96_73 in96 sn73 11140.846016
Rwneg96_74 in96 sn74 11140.846016
Rwneg96_75 in96 sn75 3183.098862
Rwneg96_76 in96 sn76 11140.846016
Rwneg96_77 in96 sn77 3183.098862
Rwneg96_78 in96 sn78 11140.846016
Rwneg96_79 in96 sn79 11140.846016
Rwneg96_80 in96 sn80 11140.846016
Rwneg96_81 in96 sn81 3183.098862
Rwneg96_82 in96 sn82 11140.846016
Rwneg96_83 in96 sn83 3183.098862
Rwneg96_84 in96 sn84 11140.846016
Rwneg96_85 in96 sn85 11140.846016
Rwneg96_86 in96 sn86 11140.846016
Rwneg96_87 in96 sn87 11140.846016
Rwneg96_88 in96 sn88 11140.846016
Rwneg96_89 in96 sn89 11140.846016
Rwneg96_90 in96 sn90 11140.846016
Rwneg96_91 in96 sn91 11140.846016
Rwneg96_92 in96 sn92 11140.846016
Rwneg96_93 in96 sn93 3183.098862
Rwneg96_94 in96 sn94 3183.098862
Rwneg96_95 in96 sn95 11140.846016
Rwneg96_96 in96 sn96 3183.098862
Rwneg96_97 in96 sn97 11140.846016
Rwneg96_98 in96 sn98 3183.098862
Rwneg96_99 in96 sn99 3183.098862
Rwneg96_100 in96 sn100 3183.098862
Rwneg97_1 in97 sn1 3183.098862
Rwneg97_2 in97 sn2 11140.846016
Rwneg97_3 in97 sn3 11140.846016
Rwneg97_4 in97 sn4 11140.846016
Rwneg97_5 in97 sn5 3183.098862
Rwneg97_6 in97 sn6 3183.098862
Rwneg97_7 in97 sn7 3183.098862
Rwneg97_8 in97 sn8 11140.846016
Rwneg97_9 in97 sn9 3183.098862
Rwneg97_10 in97 sn10 3183.098862
Rwneg97_11 in97 sn11 11140.846016
Rwneg97_12 in97 sn12 11140.846016
Rwneg97_13 in97 sn13 3183.098862
Rwneg97_14 in97 sn14 11140.846016
Rwneg97_15 in97 sn15 3183.098862
Rwneg97_16 in97 sn16 3183.098862
Rwneg97_17 in97 sn17 3183.098862
Rwneg97_18 in97 sn18 11140.846016
Rwneg97_19 in97 sn19 11140.846016
Rwneg97_20 in97 sn20 3183.098862
Rwneg97_21 in97 sn21 3183.098862
Rwneg97_22 in97 sn22 3183.098862
Rwneg97_23 in97 sn23 11140.846016
Rwneg97_24 in97 sn24 11140.846016
Rwneg97_25 in97 sn25 11140.846016
Rwneg97_26 in97 sn26 3183.098862
Rwneg97_27 in97 sn27 11140.846016
Rwneg97_28 in97 sn28 3183.098862
Rwneg97_29 in97 sn29 11140.846016
Rwneg97_30 in97 sn30 11140.846016
Rwneg97_31 in97 sn31 3183.098862
Rwneg97_32 in97 sn32 3183.098862
Rwneg97_33 in97 sn33 11140.846016
Rwneg97_34 in97 sn34 11140.846016
Rwneg97_35 in97 sn35 11140.846016
Rwneg97_36 in97 sn36 11140.846016
Rwneg97_37 in97 sn37 11140.846016
Rwneg97_38 in97 sn38 3183.098862
Rwneg97_39 in97 sn39 3183.098862
Rwneg97_40 in97 sn40 11140.846016
Rwneg97_41 in97 sn41 3183.098862
Rwneg97_42 in97 sn42 3183.098862
Rwneg97_43 in97 sn43 11140.846016
Rwneg97_44 in97 sn44 11140.846016
Rwneg97_45 in97 sn45 11140.846016
Rwneg97_46 in97 sn46 3183.098862
Rwneg97_47 in97 sn47 3183.098862
Rwneg97_48 in97 sn48 11140.846016
Rwneg97_49 in97 sn49 3183.098862
Rwneg97_50 in97 sn50 11140.846016
Rwneg97_51 in97 sn51 11140.846016
Rwneg97_52 in97 sn52 3183.098862
Rwneg97_53 in97 sn53 3183.098862
Rwneg97_54 in97 sn54 3183.098862
Rwneg97_55 in97 sn55 3183.098862
Rwneg97_56 in97 sn56 11140.846016
Rwneg97_57 in97 sn57 11140.846016
Rwneg97_58 in97 sn58 3183.098862
Rwneg97_59 in97 sn59 11140.846016
Rwneg97_60 in97 sn60 3183.098862
Rwneg97_61 in97 sn61 11140.846016
Rwneg97_62 in97 sn62 3183.098862
Rwneg97_63 in97 sn63 11140.846016
Rwneg97_64 in97 sn64 3183.098862
Rwneg97_65 in97 sn65 11140.846016
Rwneg97_66 in97 sn66 3183.098862
Rwneg97_67 in97 sn67 11140.846016
Rwneg97_68 in97 sn68 3183.098862
Rwneg97_69 in97 sn69 3183.098862
Rwneg97_70 in97 sn70 3183.098862
Rwneg97_71 in97 sn71 3183.098862
Rwneg97_72 in97 sn72 11140.846016
Rwneg97_73 in97 sn73 3183.098862
Rwneg97_74 in97 sn74 11140.846016
Rwneg97_75 in97 sn75 11140.846016
Rwneg97_76 in97 sn76 11140.846016
Rwneg97_77 in97 sn77 11140.846016
Rwneg97_78 in97 sn78 11140.846016
Rwneg97_79 in97 sn79 11140.846016
Rwneg97_80 in97 sn80 3183.098862
Rwneg97_81 in97 sn81 3183.098862
Rwneg97_82 in97 sn82 3183.098862
Rwneg97_83 in97 sn83 11140.846016
Rwneg97_84 in97 sn84 11140.846016
Rwneg97_85 in97 sn85 11140.846016
Rwneg97_86 in97 sn86 11140.846016
Rwneg97_87 in97 sn87 3183.098862
Rwneg97_88 in97 sn88 3183.098862
Rwneg97_89 in97 sn89 11140.846016
Rwneg97_90 in97 sn90 3183.098862
Rwneg97_91 in97 sn91 3183.098862
Rwneg97_92 in97 sn92 3183.098862
Rwneg97_93 in97 sn93 11140.846016
Rwneg97_94 in97 sn94 3183.098862
Rwneg97_95 in97 sn95 11140.846016
Rwneg97_96 in97 sn96 3183.098862
Rwneg97_97 in97 sn97 3183.098862
Rwneg97_98 in97 sn98 3183.098862
Rwneg97_99 in97 sn99 11140.846016
Rwneg97_100 in97 sn100 11140.846016
Rwneg98_1 in98 sn1 3183.098862
Rwneg98_2 in98 sn2 3183.098862
Rwneg98_3 in98 sn3 3183.098862
Rwneg98_4 in98 sn4 11140.846016
Rwneg98_5 in98 sn5 11140.846016
Rwneg98_6 in98 sn6 3183.098862
Rwneg98_7 in98 sn7 11140.846016
Rwneg98_8 in98 sn8 3183.098862
Rwneg98_9 in98 sn9 11140.846016
Rwneg98_10 in98 sn10 11140.846016
Rwneg98_11 in98 sn11 11140.846016
Rwneg98_12 in98 sn12 3183.098862
Rwneg98_13 in98 sn13 3183.098862
Rwneg98_14 in98 sn14 11140.846016
Rwneg98_15 in98 sn15 3183.098862
Rwneg98_16 in98 sn16 11140.846016
Rwneg98_17 in98 sn17 11140.846016
Rwneg98_18 in98 sn18 11140.846016
Rwneg98_19 in98 sn19 11140.846016
Rwneg98_20 in98 sn20 11140.846016
Rwneg98_21 in98 sn21 3183.098862
Rwneg98_22 in98 sn22 11140.846016
Rwneg98_23 in98 sn23 3183.098862
Rwneg98_24 in98 sn24 3183.098862
Rwneg98_25 in98 sn25 3183.098862
Rwneg98_26 in98 sn26 3183.098862
Rwneg98_27 in98 sn27 11140.846016
Rwneg98_28 in98 sn28 3183.098862
Rwneg98_29 in98 sn29 3183.098862
Rwneg98_30 in98 sn30 11140.846016
Rwneg98_31 in98 sn31 11140.846016
Rwneg98_32 in98 sn32 11140.846016
Rwneg98_33 in98 sn33 3183.098862
Rwneg98_34 in98 sn34 11140.846016
Rwneg98_35 in98 sn35 11140.846016
Rwneg98_36 in98 sn36 3183.098862
Rwneg98_37 in98 sn37 3183.098862
Rwneg98_38 in98 sn38 11140.846016
Rwneg98_39 in98 sn39 3183.098862
Rwneg98_40 in98 sn40 11140.846016
Rwneg98_41 in98 sn41 3183.098862
Rwneg98_42 in98 sn42 11140.846016
Rwneg98_43 in98 sn43 11140.846016
Rwneg98_44 in98 sn44 11140.846016
Rwneg98_45 in98 sn45 11140.846016
Rwneg98_46 in98 sn46 11140.846016
Rwneg98_47 in98 sn47 3183.098862
Rwneg98_48 in98 sn48 11140.846016
Rwneg98_49 in98 sn49 11140.846016
Rwneg98_50 in98 sn50 11140.846016
Rwneg98_51 in98 sn51 11140.846016
Rwneg98_52 in98 sn52 3183.098862
Rwneg98_53 in98 sn53 3183.098862
Rwneg98_54 in98 sn54 11140.846016
Rwneg98_55 in98 sn55 11140.846016
Rwneg98_56 in98 sn56 3183.098862
Rwneg98_57 in98 sn57 11140.846016
Rwneg98_58 in98 sn58 3183.098862
Rwneg98_59 in98 sn59 3183.098862
Rwneg98_60 in98 sn60 3183.098862
Rwneg98_61 in98 sn61 11140.846016
Rwneg98_62 in98 sn62 11140.846016
Rwneg98_63 in98 sn63 3183.098862
Rwneg98_64 in98 sn64 11140.846016
Rwneg98_65 in98 sn65 3183.098862
Rwneg98_66 in98 sn66 11140.846016
Rwneg98_67 in98 sn67 3183.098862
Rwneg98_68 in98 sn68 11140.846016
Rwneg98_69 in98 sn69 11140.846016
Rwneg98_70 in98 sn70 11140.846016
Rwneg98_71 in98 sn71 3183.098862
Rwneg98_72 in98 sn72 3183.098862
Rwneg98_73 in98 sn73 11140.846016
Rwneg98_74 in98 sn74 3183.098862
Rwneg98_75 in98 sn75 11140.846016
Rwneg98_76 in98 sn76 3183.098862
Rwneg98_77 in98 sn77 11140.846016
Rwneg98_78 in98 sn78 3183.098862
Rwneg98_79 in98 sn79 11140.846016
Rwneg98_80 in98 sn80 3183.098862
Rwneg98_81 in98 sn81 3183.098862
Rwneg98_82 in98 sn82 11140.846016
Rwneg98_83 in98 sn83 3183.098862
Rwneg98_84 in98 sn84 3183.098862
Rwneg98_85 in98 sn85 3183.098862
Rwneg98_86 in98 sn86 11140.846016
Rwneg98_87 in98 sn87 3183.098862
Rwneg98_88 in98 sn88 3183.098862
Rwneg98_89 in98 sn89 3183.098862
Rwneg98_90 in98 sn90 3183.098862
Rwneg98_91 in98 sn91 3183.098862
Rwneg98_92 in98 sn92 3183.098862
Rwneg98_93 in98 sn93 11140.846016
Rwneg98_94 in98 sn94 3183.098862
Rwneg98_95 in98 sn95 11140.846016
Rwneg98_96 in98 sn96 3183.098862
Rwneg98_97 in98 sn97 3183.098862
Rwneg98_98 in98 sn98 11140.846016
Rwneg98_99 in98 sn99 3183.098862
Rwneg98_100 in98 sn100 11140.846016
Rwneg99_1 in99 sn1 11140.846016
Rwneg99_2 in99 sn2 3183.098862
Rwneg99_3 in99 sn3 3183.098862
Rwneg99_4 in99 sn4 3183.098862
Rwneg99_5 in99 sn5 3183.098862
Rwneg99_6 in99 sn6 3183.098862
Rwneg99_7 in99 sn7 11140.846016
Rwneg99_8 in99 sn8 3183.098862
Rwneg99_9 in99 sn9 11140.846016
Rwneg99_10 in99 sn10 3183.098862
Rwneg99_11 in99 sn11 11140.846016
Rwneg99_12 in99 sn12 3183.098862
Rwneg99_13 in99 sn13 11140.846016
Rwneg99_14 in99 sn14 3183.098862
Rwneg99_15 in99 sn15 11140.846016
Rwneg99_16 in99 sn16 11140.846016
Rwneg99_17 in99 sn17 11140.846016
Rwneg99_18 in99 sn18 11140.846016
Rwneg99_19 in99 sn19 3183.098862
Rwneg99_20 in99 sn20 3183.098862
Rwneg99_21 in99 sn21 11140.846016
Rwneg99_22 in99 sn22 3183.098862
Rwneg99_23 in99 sn23 3183.098862
Rwneg99_24 in99 sn24 3183.098862
Rwneg99_25 in99 sn25 11140.846016
Rwneg99_26 in99 sn26 11140.846016
Rwneg99_27 in99 sn27 3183.098862
Rwneg99_28 in99 sn28 3183.098862
Rwneg99_29 in99 sn29 3183.098862
Rwneg99_30 in99 sn30 3183.098862
Rwneg99_31 in99 sn31 3183.098862
Rwneg99_32 in99 sn32 3183.098862
Rwneg99_33 in99 sn33 3183.098862
Rwneg99_34 in99 sn34 3183.098862
Rwneg99_35 in99 sn35 3183.098862
Rwneg99_36 in99 sn36 11140.846016
Rwneg99_37 in99 sn37 3183.098862
Rwneg99_38 in99 sn38 3183.098862
Rwneg99_39 in99 sn39 11140.846016
Rwneg99_40 in99 sn40 11140.846016
Rwneg99_41 in99 sn41 11140.846016
Rwneg99_42 in99 sn42 3183.098862
Rwneg99_43 in99 sn43 11140.846016
Rwneg99_44 in99 sn44 11140.846016
Rwneg99_45 in99 sn45 11140.846016
Rwneg99_46 in99 sn46 3183.098862
Rwneg99_47 in99 sn47 11140.846016
Rwneg99_48 in99 sn48 11140.846016
Rwneg99_49 in99 sn49 11140.846016
Rwneg99_50 in99 sn50 3183.098862
Rwneg99_51 in99 sn51 11140.846016
Rwneg99_52 in99 sn52 3183.098862
Rwneg99_53 in99 sn53 11140.846016
Rwneg99_54 in99 sn54 3183.098862
Rwneg99_55 in99 sn55 3183.098862
Rwneg99_56 in99 sn56 11140.846016
Rwneg99_57 in99 sn57 3183.098862
Rwneg99_58 in99 sn58 3183.098862
Rwneg99_59 in99 sn59 3183.098862
Rwneg99_60 in99 sn60 3183.098862
Rwneg99_61 in99 sn61 11140.846016
Rwneg99_62 in99 sn62 3183.098862
Rwneg99_63 in99 sn63 3183.098862
Rwneg99_64 in99 sn64 3183.098862
Rwneg99_65 in99 sn65 11140.846016
Rwneg99_66 in99 sn66 3183.098862
Rwneg99_67 in99 sn67 3183.098862
Rwneg99_68 in99 sn68 11140.846016
Rwneg99_69 in99 sn69 3183.098862
Rwneg99_70 in99 sn70 3183.098862
Rwneg99_71 in99 sn71 11140.846016
Rwneg99_72 in99 sn72 3183.098862
Rwneg99_73 in99 sn73 3183.098862
Rwneg99_74 in99 sn74 11140.846016
Rwneg99_75 in99 sn75 11140.846016
Rwneg99_76 in99 sn76 11140.846016
Rwneg99_77 in99 sn77 3183.098862
Rwneg99_78 in99 sn78 11140.846016
Rwneg99_79 in99 sn79 11140.846016
Rwneg99_80 in99 sn80 11140.846016
Rwneg99_81 in99 sn81 11140.846016
Rwneg99_82 in99 sn82 11140.846016
Rwneg99_83 in99 sn83 11140.846016
Rwneg99_84 in99 sn84 11140.846016
Rwneg99_85 in99 sn85 3183.098862
Rwneg99_86 in99 sn86 3183.098862
Rwneg99_87 in99 sn87 11140.846016
Rwneg99_88 in99 sn88 3183.098862
Rwneg99_89 in99 sn89 11140.846016
Rwneg99_90 in99 sn90 3183.098862
Rwneg99_91 in99 sn91 11140.846016
Rwneg99_92 in99 sn92 11140.846016
Rwneg99_93 in99 sn93 3183.098862
Rwneg99_94 in99 sn94 3183.098862
Rwneg99_95 in99 sn95 3183.098862
Rwneg99_96 in99 sn96 11140.846016
Rwneg99_97 in99 sn97 3183.098862
Rwneg99_98 in99 sn98 11140.846016
Rwneg99_99 in99 sn99 3183.098862
Rwneg99_100 in99 sn100 3183.098862
Rwneg100_1 in100 sn1 3183.098862
Rwneg100_2 in100 sn2 3183.098862
Rwneg100_3 in100 sn3 3183.098862
Rwneg100_4 in100 sn4 3183.098862
Rwneg100_5 in100 sn5 3183.098862
Rwneg100_6 in100 sn6 3183.098862
Rwneg100_7 in100 sn7 11140.846016
Rwneg100_8 in100 sn8 3183.098862
Rwneg100_9 in100 sn9 3183.098862
Rwneg100_10 in100 sn10 11140.846016
Rwneg100_11 in100 sn11 11140.846016
Rwneg100_12 in100 sn12 11140.846016
Rwneg100_13 in100 sn13 11140.846016
Rwneg100_14 in100 sn14 3183.098862
Rwneg100_15 in100 sn15 3183.098862
Rwneg100_16 in100 sn16 3183.098862
Rwneg100_17 in100 sn17 11140.846016
Rwneg100_18 in100 sn18 11140.846016
Rwneg100_19 in100 sn19 11140.846016
Rwneg100_20 in100 sn20 11140.846016
Rwneg100_21 in100 sn21 3183.098862
Rwneg100_22 in100 sn22 11140.846016
Rwneg100_23 in100 sn23 11140.846016
Rwneg100_24 in100 sn24 11140.846016
Rwneg100_25 in100 sn25 3183.098862
Rwneg100_26 in100 sn26 3183.098862
Rwneg100_27 in100 sn27 11140.846016
Rwneg100_28 in100 sn28 11140.846016
Rwneg100_29 in100 sn29 11140.846016
Rwneg100_30 in100 sn30 11140.846016
Rwneg100_31 in100 sn31 3183.098862
Rwneg100_32 in100 sn32 11140.846016
Rwneg100_33 in100 sn33 11140.846016
Rwneg100_34 in100 sn34 11140.846016
Rwneg100_35 in100 sn35 11140.846016
Rwneg100_36 in100 sn36 11140.846016
Rwneg100_37 in100 sn37 3183.098862
Rwneg100_38 in100 sn38 11140.846016
Rwneg100_39 in100 sn39 11140.846016
Rwneg100_40 in100 sn40 11140.846016
Rwneg100_41 in100 sn41 11140.846016
Rwneg100_42 in100 sn42 3183.098862
Rwneg100_43 in100 sn43 3183.098862
Rwneg100_44 in100 sn44 11140.846016
Rwneg100_45 in100 sn45 11140.846016
Rwneg100_46 in100 sn46 3183.098862
Rwneg100_47 in100 sn47 3183.098862
Rwneg100_48 in100 sn48 3183.098862
Rwneg100_49 in100 sn49 11140.846016
Rwneg100_50 in100 sn50 11140.846016
Rwneg100_51 in100 sn51 3183.098862
Rwneg100_52 in100 sn52 3183.098862
Rwneg100_53 in100 sn53 11140.846016
Rwneg100_54 in100 sn54 3183.098862
Rwneg100_55 in100 sn55 11140.846016
Rwneg100_56 in100 sn56 3183.098862
Rwneg100_57 in100 sn57 11140.846016
Rwneg100_58 in100 sn58 3183.098862
Rwneg100_59 in100 sn59 3183.098862
Rwneg100_60 in100 sn60 11140.846016
Rwneg100_61 in100 sn61 11140.846016
Rwneg100_62 in100 sn62 11140.846016
Rwneg100_63 in100 sn63 3183.098862
Rwneg100_64 in100 sn64 3183.098862
Rwneg100_65 in100 sn65 11140.846016
Rwneg100_66 in100 sn66 3183.098862
Rwneg100_67 in100 sn67 11140.846016
Rwneg100_68 in100 sn68 3183.098862
Rwneg100_69 in100 sn69 3183.098862
Rwneg100_70 in100 sn70 3183.098862
Rwneg100_71 in100 sn71 11140.846016
Rwneg100_72 in100 sn72 11140.846016
Rwneg100_73 in100 sn73 11140.846016
Rwneg100_74 in100 sn74 11140.846016
Rwneg100_75 in100 sn75 11140.846016
Rwneg100_76 in100 sn76 11140.846016
Rwneg100_77 in100 sn77 11140.846016
Rwneg100_78 in100 sn78 11140.846016
Rwneg100_79 in100 sn79 3183.098862
Rwneg100_80 in100 sn80 3183.098862
Rwneg100_81 in100 sn81 3183.098862
Rwneg100_82 in100 sn82 11140.846016
Rwneg100_83 in100 sn83 11140.846016
Rwneg100_84 in100 sn84 11140.846016
Rwneg100_85 in100 sn85 11140.846016
Rwneg100_86 in100 sn86 3183.098862
Rwneg100_87 in100 sn87 11140.846016
Rwneg100_88 in100 sn88 3183.098862
Rwneg100_89 in100 sn89 3183.098862
Rwneg100_90 in100 sn90 3183.098862
Rwneg100_91 in100 sn91 3183.098862
Rwneg100_92 in100 sn92 11140.846016
Rwneg100_93 in100 sn93 3183.098862
Rwneg100_94 in100 sn94 11140.846016
Rwneg100_95 in100 sn95 11140.846016
Rwneg100_96 in100 sn96 3183.098862
Rwneg100_97 in100 sn97 11140.846016
Rwneg100_98 in100 sn98 11140.846016
Rwneg100_99 in100 sn99 3183.098862
Rwneg100_100 in100 sn100 3183.098862
Rwneg101_1 in101 sn1 3183.098862
Rwneg101_2 in101 sn2 11140.846016
Rwneg101_3 in101 sn3 11140.846016
Rwneg101_4 in101 sn4 3183.098862
Rwneg101_5 in101 sn5 11140.846016
Rwneg101_6 in101 sn6 3183.098862
Rwneg101_7 in101 sn7 3183.098862
Rwneg101_8 in101 sn8 11140.846016
Rwneg101_9 in101 sn9 3183.098862
Rwneg101_10 in101 sn10 11140.846016
Rwneg101_11 in101 sn11 3183.098862
Rwneg101_12 in101 sn12 3183.098862
Rwneg101_13 in101 sn13 3183.098862
Rwneg101_14 in101 sn14 11140.846016
Rwneg101_15 in101 sn15 3183.098862
Rwneg101_16 in101 sn16 11140.846016
Rwneg101_17 in101 sn17 11140.846016
Rwneg101_18 in101 sn18 11140.846016
Rwneg101_19 in101 sn19 11140.846016
Rwneg101_20 in101 sn20 11140.846016
Rwneg101_21 in101 sn21 11140.846016
Rwneg101_22 in101 sn22 11140.846016
Rwneg101_23 in101 sn23 3183.098862
Rwneg101_24 in101 sn24 11140.846016
Rwneg101_25 in101 sn25 3183.098862
Rwneg101_26 in101 sn26 11140.846016
Rwneg101_27 in101 sn27 11140.846016
Rwneg101_28 in101 sn28 3183.098862
Rwneg101_29 in101 sn29 11140.846016
Rwneg101_30 in101 sn30 11140.846016
Rwneg101_31 in101 sn31 3183.098862
Rwneg101_32 in101 sn32 11140.846016
Rwneg101_33 in101 sn33 3183.098862
Rwneg101_34 in101 sn34 3183.098862
Rwneg101_35 in101 sn35 11140.846016
Rwneg101_36 in101 sn36 11140.846016
Rwneg101_37 in101 sn37 11140.846016
Rwneg101_38 in101 sn38 3183.098862
Rwneg101_39 in101 sn39 11140.846016
Rwneg101_40 in101 sn40 11140.846016
Rwneg101_41 in101 sn41 3183.098862
Rwneg101_42 in101 sn42 11140.846016
Rwneg101_43 in101 sn43 11140.846016
Rwneg101_44 in101 sn44 11140.846016
Rwneg101_45 in101 sn45 3183.098862
Rwneg101_46 in101 sn46 11140.846016
Rwneg101_47 in101 sn47 11140.846016
Rwneg101_48 in101 sn48 11140.846016
Rwneg101_49 in101 sn49 11140.846016
Rwneg101_50 in101 sn50 3183.098862
Rwneg101_51 in101 sn51 11140.846016
Rwneg101_52 in101 sn52 11140.846016
Rwneg101_53 in101 sn53 3183.098862
Rwneg101_54 in101 sn54 11140.846016
Rwneg101_55 in101 sn55 11140.846016
Rwneg101_56 in101 sn56 3183.098862
Rwneg101_57 in101 sn57 3183.098862
Rwneg101_58 in101 sn58 11140.846016
Rwneg101_59 in101 sn59 11140.846016
Rwneg101_60 in101 sn60 3183.098862
Rwneg101_61 in101 sn61 3183.098862
Rwneg101_62 in101 sn62 11140.846016
Rwneg101_63 in101 sn63 3183.098862
Rwneg101_64 in101 sn64 11140.846016
Rwneg101_65 in101 sn65 3183.098862
Rwneg101_66 in101 sn66 3183.098862
Rwneg101_67 in101 sn67 11140.846016
Rwneg101_68 in101 sn68 11140.846016
Rwneg101_69 in101 sn69 3183.098862
Rwneg101_70 in101 sn70 11140.846016
Rwneg101_71 in101 sn71 11140.846016
Rwneg101_72 in101 sn72 3183.098862
Rwneg101_73 in101 sn73 3183.098862
Rwneg101_74 in101 sn74 11140.846016
Rwneg101_75 in101 sn75 11140.846016
Rwneg101_76 in101 sn76 11140.846016
Rwneg101_77 in101 sn77 3183.098862
Rwneg101_78 in101 sn78 3183.098862
Rwneg101_79 in101 sn79 3183.098862
Rwneg101_80 in101 sn80 11140.846016
Rwneg101_81 in101 sn81 3183.098862
Rwneg101_82 in101 sn82 3183.098862
Rwneg101_83 in101 sn83 11140.846016
Rwneg101_84 in101 sn84 11140.846016
Rwneg101_85 in101 sn85 11140.846016
Rwneg101_86 in101 sn86 11140.846016
Rwneg101_87 in101 sn87 11140.846016
Rwneg101_88 in101 sn88 11140.846016
Rwneg101_89 in101 sn89 11140.846016
Rwneg101_90 in101 sn90 3183.098862
Rwneg101_91 in101 sn91 11140.846016
Rwneg101_92 in101 sn92 3183.098862
Rwneg101_93 in101 sn93 3183.098862
Rwneg101_94 in101 sn94 11140.846016
Rwneg101_95 in101 sn95 3183.098862
Rwneg101_96 in101 sn96 11140.846016
Rwneg101_97 in101 sn97 3183.098862
Rwneg101_98 in101 sn98 3183.098862
Rwneg101_99 in101 sn99 11140.846016
Rwneg101_100 in101 sn100 3183.098862
Rwneg102_1 in102 sn1 11140.846016
Rwneg102_2 in102 sn2 11140.846016
Rwneg102_3 in102 sn3 3183.098862
Rwneg102_4 in102 sn4 3183.098862
Rwneg102_5 in102 sn5 3183.098862
Rwneg102_6 in102 sn6 11140.846016
Rwneg102_7 in102 sn7 11140.846016
Rwneg102_8 in102 sn8 11140.846016
Rwneg102_9 in102 sn9 3183.098862
Rwneg102_10 in102 sn10 3183.098862
Rwneg102_11 in102 sn11 3183.098862
Rwneg102_12 in102 sn12 11140.846016
Rwneg102_13 in102 sn13 11140.846016
Rwneg102_14 in102 sn14 3183.098862
Rwneg102_15 in102 sn15 11140.846016
Rwneg102_16 in102 sn16 3183.098862
Rwneg102_17 in102 sn17 3183.098862
Rwneg102_18 in102 sn18 3183.098862
Rwneg102_19 in102 sn19 3183.098862
Rwneg102_20 in102 sn20 3183.098862
Rwneg102_21 in102 sn21 3183.098862
Rwneg102_22 in102 sn22 3183.098862
Rwneg102_23 in102 sn23 11140.846016
Rwneg102_24 in102 sn24 11140.846016
Rwneg102_25 in102 sn25 11140.846016
Rwneg102_26 in102 sn26 11140.846016
Rwneg102_27 in102 sn27 11140.846016
Rwneg102_28 in102 sn28 11140.846016
Rwneg102_29 in102 sn29 11140.846016
Rwneg102_30 in102 sn30 11140.846016
Rwneg102_31 in102 sn31 11140.846016
Rwneg102_32 in102 sn32 11140.846016
Rwneg102_33 in102 sn33 11140.846016
Rwneg102_34 in102 sn34 11140.846016
Rwneg102_35 in102 sn35 3183.098862
Rwneg102_36 in102 sn36 11140.846016
Rwneg102_37 in102 sn37 3183.098862
Rwneg102_38 in102 sn38 11140.846016
Rwneg102_39 in102 sn39 3183.098862
Rwneg102_40 in102 sn40 11140.846016
Rwneg102_41 in102 sn41 3183.098862
Rwneg102_42 in102 sn42 3183.098862
Rwneg102_43 in102 sn43 11140.846016
Rwneg102_44 in102 sn44 3183.098862
Rwneg102_45 in102 sn45 11140.846016
Rwneg102_46 in102 sn46 3183.098862
Rwneg102_47 in102 sn47 11140.846016
Rwneg102_48 in102 sn48 3183.098862
Rwneg102_49 in102 sn49 3183.098862
Rwneg102_50 in102 sn50 3183.098862
Rwneg102_51 in102 sn51 11140.846016
Rwneg102_52 in102 sn52 3183.098862
Rwneg102_53 in102 sn53 3183.098862
Rwneg102_54 in102 sn54 11140.846016
Rwneg102_55 in102 sn55 3183.098862
Rwneg102_56 in102 sn56 11140.846016
Rwneg102_57 in102 sn57 11140.846016
Rwneg102_58 in102 sn58 3183.098862
Rwneg102_59 in102 sn59 11140.846016
Rwneg102_60 in102 sn60 3183.098862
Rwneg102_61 in102 sn61 3183.098862
Rwneg102_62 in102 sn62 3183.098862
Rwneg102_63 in102 sn63 11140.846016
Rwneg102_64 in102 sn64 11140.846016
Rwneg102_65 in102 sn65 11140.846016
Rwneg102_66 in102 sn66 3183.098862
Rwneg102_67 in102 sn67 11140.846016
Rwneg102_68 in102 sn68 11140.846016
Rwneg102_69 in102 sn69 3183.098862
Rwneg102_70 in102 sn70 3183.098862
Rwneg102_71 in102 sn71 3183.098862
Rwneg102_72 in102 sn72 3183.098862
Rwneg102_73 in102 sn73 3183.098862
Rwneg102_74 in102 sn74 11140.846016
Rwneg102_75 in102 sn75 11140.846016
Rwneg102_76 in102 sn76 3183.098862
Rwneg102_77 in102 sn77 11140.846016
Rwneg102_78 in102 sn78 3183.098862
Rwneg102_79 in102 sn79 11140.846016
Rwneg102_80 in102 sn80 11140.846016
Rwneg102_81 in102 sn81 11140.846016
Rwneg102_82 in102 sn82 11140.846016
Rwneg102_83 in102 sn83 11140.846016
Rwneg102_84 in102 sn84 11140.846016
Rwneg102_85 in102 sn85 11140.846016
Rwneg102_86 in102 sn86 11140.846016
Rwneg102_87 in102 sn87 3183.098862
Rwneg102_88 in102 sn88 3183.098862
Rwneg102_89 in102 sn89 3183.098862
Rwneg102_90 in102 sn90 3183.098862
Rwneg102_91 in102 sn91 11140.846016
Rwneg102_92 in102 sn92 3183.098862
Rwneg102_93 in102 sn93 3183.098862
Rwneg102_94 in102 sn94 11140.846016
Rwneg102_95 in102 sn95 11140.846016
Rwneg102_96 in102 sn96 11140.846016
Rwneg102_97 in102 sn97 11140.846016
Rwneg102_98 in102 sn98 3183.098862
Rwneg102_99 in102 sn99 3183.098862
Rwneg102_100 in102 sn100 11140.846016
Rwneg103_1 in103 sn1 3183.098862
Rwneg103_2 in103 sn2 11140.846016
Rwneg103_3 in103 sn3 3183.098862
Rwneg103_4 in103 sn4 3183.098862
Rwneg103_5 in103 sn5 3183.098862
Rwneg103_6 in103 sn6 3183.098862
Rwneg103_7 in103 sn7 11140.846016
Rwneg103_8 in103 sn8 3183.098862
Rwneg103_9 in103 sn9 11140.846016
Rwneg103_10 in103 sn10 3183.098862
Rwneg103_11 in103 sn11 11140.846016
Rwneg103_12 in103 sn12 11140.846016
Rwneg103_13 in103 sn13 3183.098862
Rwneg103_14 in103 sn14 11140.846016
Rwneg103_15 in103 sn15 3183.098862
Rwneg103_16 in103 sn16 3183.098862
Rwneg103_17 in103 sn17 3183.098862
Rwneg103_18 in103 sn18 11140.846016
Rwneg103_19 in103 sn19 3183.098862
Rwneg103_20 in103 sn20 3183.098862
Rwneg103_21 in103 sn21 11140.846016
Rwneg103_22 in103 sn22 3183.098862
Rwneg103_23 in103 sn23 11140.846016
Rwneg103_24 in103 sn24 3183.098862
Rwneg103_25 in103 sn25 3183.098862
Rwneg103_26 in103 sn26 11140.846016
Rwneg103_27 in103 sn27 3183.098862
Rwneg103_28 in103 sn28 11140.846016
Rwneg103_29 in103 sn29 3183.098862
Rwneg103_30 in103 sn30 11140.846016
Rwneg103_31 in103 sn31 11140.846016
Rwneg103_32 in103 sn32 3183.098862
Rwneg103_33 in103 sn33 11140.846016
Rwneg103_34 in103 sn34 3183.098862
Rwneg103_35 in103 sn35 3183.098862
Rwneg103_36 in103 sn36 11140.846016
Rwneg103_37 in103 sn37 11140.846016
Rwneg103_38 in103 sn38 3183.098862
Rwneg103_39 in103 sn39 3183.098862
Rwneg103_40 in103 sn40 3183.098862
Rwneg103_41 in103 sn41 3183.098862
Rwneg103_42 in103 sn42 11140.846016
Rwneg103_43 in103 sn43 3183.098862
Rwneg103_44 in103 sn44 11140.846016
Rwneg103_45 in103 sn45 11140.846016
Rwneg103_46 in103 sn46 11140.846016
Rwneg103_47 in103 sn47 3183.098862
Rwneg103_48 in103 sn48 11140.846016
Rwneg103_49 in103 sn49 3183.098862
Rwneg103_50 in103 sn50 11140.846016
Rwneg103_51 in103 sn51 3183.098862
Rwneg103_52 in103 sn52 3183.098862
Rwneg103_53 in103 sn53 11140.846016
Rwneg103_54 in103 sn54 3183.098862
Rwneg103_55 in103 sn55 11140.846016
Rwneg103_56 in103 sn56 3183.098862
Rwneg103_57 in103 sn57 11140.846016
Rwneg103_58 in103 sn58 3183.098862
Rwneg103_59 in103 sn59 11140.846016
Rwneg103_60 in103 sn60 3183.098862
Rwneg103_61 in103 sn61 11140.846016
Rwneg103_62 in103 sn62 3183.098862
Rwneg103_63 in103 sn63 3183.098862
Rwneg103_64 in103 sn64 3183.098862
Rwneg103_65 in103 sn65 3183.098862
Rwneg103_66 in103 sn66 11140.846016
Rwneg103_67 in103 sn67 11140.846016
Rwneg103_68 in103 sn68 3183.098862
Rwneg103_69 in103 sn69 11140.846016
Rwneg103_70 in103 sn70 3183.098862
Rwneg103_71 in103 sn71 11140.846016
Rwneg103_72 in103 sn72 11140.846016
Rwneg103_73 in103 sn73 11140.846016
Rwneg103_74 in103 sn74 3183.098862
Rwneg103_75 in103 sn75 3183.098862
Rwneg103_76 in103 sn76 3183.098862
Rwneg103_77 in103 sn77 11140.846016
Rwneg103_78 in103 sn78 3183.098862
Rwneg103_79 in103 sn79 11140.846016
Rwneg103_80 in103 sn80 3183.098862
Rwneg103_81 in103 sn81 3183.098862
Rwneg103_82 in103 sn82 11140.846016
Rwneg103_83 in103 sn83 3183.098862
Rwneg103_84 in103 sn84 11140.846016
Rwneg103_85 in103 sn85 3183.098862
Rwneg103_86 in103 sn86 3183.098862
Rwneg103_87 in103 sn87 3183.098862
Rwneg103_88 in103 sn88 11140.846016
Rwneg103_89 in103 sn89 11140.846016
Rwneg103_90 in103 sn90 11140.846016
Rwneg103_91 in103 sn91 3183.098862
Rwneg103_92 in103 sn92 3183.098862
Rwneg103_93 in103 sn93 3183.098862
Rwneg103_94 in103 sn94 3183.098862
Rwneg103_95 in103 sn95 11140.846016
Rwneg103_96 in103 sn96 3183.098862
Rwneg103_97 in103 sn97 3183.098862
Rwneg103_98 in103 sn98 3183.098862
Rwneg103_99 in103 sn99 11140.846016
Rwneg103_100 in103 sn100 11140.846016
Rwneg104_1 in104 sn1 3183.098862
Rwneg104_2 in104 sn2 3183.098862
Rwneg104_3 in104 sn3 11140.846016
Rwneg104_4 in104 sn4 11140.846016
Rwneg104_5 in104 sn5 3183.098862
Rwneg104_6 in104 sn6 3183.098862
Rwneg104_7 in104 sn7 3183.098862
Rwneg104_8 in104 sn8 11140.846016
Rwneg104_9 in104 sn9 11140.846016
Rwneg104_10 in104 sn10 11140.846016
Rwneg104_11 in104 sn11 3183.098862
Rwneg104_12 in104 sn12 11140.846016
Rwneg104_13 in104 sn13 3183.098862
Rwneg104_14 in104 sn14 11140.846016
Rwneg104_15 in104 sn15 3183.098862
Rwneg104_16 in104 sn16 3183.098862
Rwneg104_17 in104 sn17 3183.098862
Rwneg104_18 in104 sn18 3183.098862
Rwneg104_19 in104 sn19 11140.846016
Rwneg104_20 in104 sn20 3183.098862
Rwneg104_21 in104 sn21 3183.098862
Rwneg104_22 in104 sn22 3183.098862
Rwneg104_23 in104 sn23 11140.846016
Rwneg104_24 in104 sn24 3183.098862
Rwneg104_25 in104 sn25 3183.098862
Rwneg104_26 in104 sn26 11140.846016
Rwneg104_27 in104 sn27 11140.846016
Rwneg104_28 in104 sn28 11140.846016
Rwneg104_29 in104 sn29 11140.846016
Rwneg104_30 in104 sn30 3183.098862
Rwneg104_31 in104 sn31 3183.098862
Rwneg104_32 in104 sn32 3183.098862
Rwneg104_33 in104 sn33 3183.098862
Rwneg104_34 in104 sn34 3183.098862
Rwneg104_35 in104 sn35 3183.098862
Rwneg104_36 in104 sn36 3183.098862
Rwneg104_37 in104 sn37 11140.846016
Rwneg104_38 in104 sn38 3183.098862
Rwneg104_39 in104 sn39 3183.098862
Rwneg104_40 in104 sn40 3183.098862
Rwneg104_41 in104 sn41 11140.846016
Rwneg104_42 in104 sn42 3183.098862
Rwneg104_43 in104 sn43 11140.846016
Rwneg104_44 in104 sn44 11140.846016
Rwneg104_45 in104 sn45 3183.098862
Rwneg104_46 in104 sn46 11140.846016
Rwneg104_47 in104 sn47 3183.098862
Rwneg104_48 in104 sn48 11140.846016
Rwneg104_49 in104 sn49 3183.098862
Rwneg104_50 in104 sn50 3183.098862
Rwneg104_51 in104 sn51 11140.846016
Rwneg104_52 in104 sn52 11140.846016
Rwneg104_53 in104 sn53 3183.098862
Rwneg104_54 in104 sn54 3183.098862
Rwneg104_55 in104 sn55 3183.098862
Rwneg104_56 in104 sn56 11140.846016
Rwneg104_57 in104 sn57 11140.846016
Rwneg104_58 in104 sn58 3183.098862
Rwneg104_59 in104 sn59 3183.098862
Rwneg104_60 in104 sn60 11140.846016
Rwneg104_61 in104 sn61 3183.098862
Rwneg104_62 in104 sn62 11140.846016
Rwneg104_63 in104 sn63 11140.846016
Rwneg104_64 in104 sn64 11140.846016
Rwneg104_65 in104 sn65 3183.098862
Rwneg104_66 in104 sn66 3183.098862
Rwneg104_67 in104 sn67 3183.098862
Rwneg104_68 in104 sn68 11140.846016
Rwneg104_69 in104 sn69 3183.098862
Rwneg104_70 in104 sn70 11140.846016
Rwneg104_71 in104 sn71 3183.098862
Rwneg104_72 in104 sn72 11140.846016
Rwneg104_73 in104 sn73 3183.098862
Rwneg104_74 in104 sn74 3183.098862
Rwneg104_75 in104 sn75 11140.846016
Rwneg104_76 in104 sn76 11140.846016
Rwneg104_77 in104 sn77 3183.098862
Rwneg104_78 in104 sn78 11140.846016
Rwneg104_79 in104 sn79 3183.098862
Rwneg104_80 in104 sn80 11140.846016
Rwneg104_81 in104 sn81 11140.846016
Rwneg104_82 in104 sn82 3183.098862
Rwneg104_83 in104 sn83 11140.846016
Rwneg104_84 in104 sn84 3183.098862
Rwneg104_85 in104 sn85 3183.098862
Rwneg104_86 in104 sn86 11140.846016
Rwneg104_87 in104 sn87 11140.846016
Rwneg104_88 in104 sn88 3183.098862
Rwneg104_89 in104 sn89 11140.846016
Rwneg104_90 in104 sn90 3183.098862
Rwneg104_91 in104 sn91 3183.098862
Rwneg104_92 in104 sn92 11140.846016
Rwneg104_93 in104 sn93 3183.098862
Rwneg104_94 in104 sn94 11140.846016
Rwneg104_95 in104 sn95 11140.846016
Rwneg104_96 in104 sn96 3183.098862
Rwneg104_97 in104 sn97 3183.098862
Rwneg104_98 in104 sn98 11140.846016
Rwneg104_99 in104 sn99 11140.846016
Rwneg104_100 in104 sn100 11140.846016
Rwneg105_1 in105 sn1 3183.098862
Rwneg105_2 in105 sn2 11140.846016
Rwneg105_3 in105 sn3 11140.846016
Rwneg105_4 in105 sn4 3183.098862
Rwneg105_5 in105 sn5 11140.846016
Rwneg105_6 in105 sn6 3183.098862
Rwneg105_7 in105 sn7 11140.846016
Rwneg105_8 in105 sn8 3183.098862
Rwneg105_9 in105 sn9 3183.098862
Rwneg105_10 in105 sn10 11140.846016
Rwneg105_11 in105 sn11 3183.098862
Rwneg105_12 in105 sn12 11140.846016
Rwneg105_13 in105 sn13 11140.846016
Rwneg105_14 in105 sn14 11140.846016
Rwneg105_15 in105 sn15 11140.846016
Rwneg105_16 in105 sn16 3183.098862
Rwneg105_17 in105 sn17 3183.098862
Rwneg105_18 in105 sn18 11140.846016
Rwneg105_19 in105 sn19 11140.846016
Rwneg105_20 in105 sn20 3183.098862
Rwneg105_21 in105 sn21 3183.098862
Rwneg105_22 in105 sn22 3183.098862
Rwneg105_23 in105 sn23 3183.098862
Rwneg105_24 in105 sn24 3183.098862
Rwneg105_25 in105 sn25 3183.098862
Rwneg105_26 in105 sn26 11140.846016
Rwneg105_27 in105 sn27 3183.098862
Rwneg105_28 in105 sn28 3183.098862
Rwneg105_29 in105 sn29 11140.846016
Rwneg105_30 in105 sn30 11140.846016
Rwneg105_31 in105 sn31 11140.846016
Rwneg105_32 in105 sn32 3183.098862
Rwneg105_33 in105 sn33 3183.098862
Rwneg105_34 in105 sn34 3183.098862
Rwneg105_35 in105 sn35 11140.846016
Rwneg105_36 in105 sn36 3183.098862
Rwneg105_37 in105 sn37 3183.098862
Rwneg105_38 in105 sn38 11140.846016
Rwneg105_39 in105 sn39 3183.098862
Rwneg105_40 in105 sn40 11140.846016
Rwneg105_41 in105 sn41 3183.098862
Rwneg105_42 in105 sn42 11140.846016
Rwneg105_43 in105 sn43 3183.098862
Rwneg105_44 in105 sn44 11140.846016
Rwneg105_45 in105 sn45 3183.098862
Rwneg105_46 in105 sn46 11140.846016
Rwneg105_47 in105 sn47 3183.098862
Rwneg105_48 in105 sn48 11140.846016
Rwneg105_49 in105 sn49 3183.098862
Rwneg105_50 in105 sn50 11140.846016
Rwneg105_51 in105 sn51 11140.846016
Rwneg105_52 in105 sn52 11140.846016
Rwneg105_53 in105 sn53 3183.098862
Rwneg105_54 in105 sn54 3183.098862
Rwneg105_55 in105 sn55 11140.846016
Rwneg105_56 in105 sn56 11140.846016
Rwneg105_57 in105 sn57 11140.846016
Rwneg105_58 in105 sn58 11140.846016
Rwneg105_59 in105 sn59 11140.846016
Rwneg105_60 in105 sn60 11140.846016
Rwneg105_61 in105 sn61 11140.846016
Rwneg105_62 in105 sn62 3183.098862
Rwneg105_63 in105 sn63 11140.846016
Rwneg105_64 in105 sn64 3183.098862
Rwneg105_65 in105 sn65 3183.098862
Rwneg105_66 in105 sn66 3183.098862
Rwneg105_67 in105 sn67 11140.846016
Rwneg105_68 in105 sn68 3183.098862
Rwneg105_69 in105 sn69 11140.846016
Rwneg105_70 in105 sn70 3183.098862
Rwneg105_71 in105 sn71 3183.098862
Rwneg105_72 in105 sn72 3183.098862
Rwneg105_73 in105 sn73 11140.846016
Rwneg105_74 in105 sn74 11140.846016
Rwneg105_75 in105 sn75 11140.846016
Rwneg105_76 in105 sn76 11140.846016
Rwneg105_77 in105 sn77 3183.098862
Rwneg105_78 in105 sn78 11140.846016
Rwneg105_79 in105 sn79 11140.846016
Rwneg105_80 in105 sn80 3183.098862
Rwneg105_81 in105 sn81 3183.098862
Rwneg105_82 in105 sn82 3183.098862
Rwneg105_83 in105 sn83 11140.846016
Rwneg105_84 in105 sn84 11140.846016
Rwneg105_85 in105 sn85 11140.846016
Rwneg105_86 in105 sn86 11140.846016
Rwneg105_87 in105 sn87 3183.098862
Rwneg105_88 in105 sn88 11140.846016
Rwneg105_89 in105 sn89 11140.846016
Rwneg105_90 in105 sn90 11140.846016
Rwneg105_91 in105 sn91 3183.098862
Rwneg105_92 in105 sn92 3183.098862
Rwneg105_93 in105 sn93 3183.098862
Rwneg105_94 in105 sn94 11140.846016
Rwneg105_95 in105 sn95 3183.098862
Rwneg105_96 in105 sn96 11140.846016
Rwneg105_97 in105 sn97 3183.098862
Rwneg105_98 in105 sn98 3183.098862
Rwneg105_99 in105 sn99 3183.098862
Rwneg105_100 in105 sn100 3183.098862
Rwneg106_1 in106 sn1 11140.846016
Rwneg106_2 in106 sn2 3183.098862
Rwneg106_3 in106 sn3 11140.846016
Rwneg106_4 in106 sn4 11140.846016
Rwneg106_5 in106 sn5 3183.098862
Rwneg106_6 in106 sn6 11140.846016
Rwneg106_7 in106 sn7 11140.846016
Rwneg106_8 in106 sn8 11140.846016
Rwneg106_9 in106 sn9 3183.098862
Rwneg106_10 in106 sn10 3183.098862
Rwneg106_11 in106 sn11 11140.846016
Rwneg106_12 in106 sn12 11140.846016
Rwneg106_13 in106 sn13 3183.098862
Rwneg106_14 in106 sn14 3183.098862
Rwneg106_15 in106 sn15 11140.846016
Rwneg106_16 in106 sn16 11140.846016
Rwneg106_17 in106 sn17 11140.846016
Rwneg106_18 in106 sn18 3183.098862
Rwneg106_19 in106 sn19 3183.098862
Rwneg106_20 in106 sn20 3183.098862
Rwneg106_21 in106 sn21 3183.098862
Rwneg106_22 in106 sn22 11140.846016
Rwneg106_23 in106 sn23 11140.846016
Rwneg106_24 in106 sn24 11140.846016
Rwneg106_25 in106 sn25 3183.098862
Rwneg106_26 in106 sn26 3183.098862
Rwneg106_27 in106 sn27 3183.098862
Rwneg106_28 in106 sn28 11140.846016
Rwneg106_29 in106 sn29 11140.846016
Rwneg106_30 in106 sn30 3183.098862
Rwneg106_31 in106 sn31 11140.846016
Rwneg106_32 in106 sn32 3183.098862
Rwneg106_33 in106 sn33 3183.098862
Rwneg106_34 in106 sn34 11140.846016
Rwneg106_35 in106 sn35 11140.846016
Rwneg106_36 in106 sn36 11140.846016
Rwneg106_37 in106 sn37 3183.098862
Rwneg106_38 in106 sn38 11140.846016
Rwneg106_39 in106 sn39 11140.846016
Rwneg106_40 in106 sn40 11140.846016
Rwneg106_41 in106 sn41 3183.098862
Rwneg106_42 in106 sn42 3183.098862
Rwneg106_43 in106 sn43 3183.098862
Rwneg106_44 in106 sn44 11140.846016
Rwneg106_45 in106 sn45 3183.098862
Rwneg106_46 in106 sn46 3183.098862
Rwneg106_47 in106 sn47 11140.846016
Rwneg106_48 in106 sn48 3183.098862
Rwneg106_49 in106 sn49 11140.846016
Rwneg106_50 in106 sn50 3183.098862
Rwneg106_51 in106 sn51 3183.098862
Rwneg106_52 in106 sn52 11140.846016
Rwneg106_53 in106 sn53 11140.846016
Rwneg106_54 in106 sn54 11140.846016
Rwneg106_55 in106 sn55 11140.846016
Rwneg106_56 in106 sn56 11140.846016
Rwneg106_57 in106 sn57 3183.098862
Rwneg106_58 in106 sn58 3183.098862
Rwneg106_59 in106 sn59 3183.098862
Rwneg106_60 in106 sn60 11140.846016
Rwneg106_61 in106 sn61 11140.846016
Rwneg106_62 in106 sn62 3183.098862
Rwneg106_63 in106 sn63 11140.846016
Rwneg106_64 in106 sn64 11140.846016
Rwneg106_65 in106 sn65 3183.098862
Rwneg106_66 in106 sn66 11140.846016
Rwneg106_67 in106 sn67 3183.098862
Rwneg106_68 in106 sn68 11140.846016
Rwneg106_69 in106 sn69 11140.846016
Rwneg106_70 in106 sn70 3183.098862
Rwneg106_71 in106 sn71 11140.846016
Rwneg106_72 in106 sn72 3183.098862
Rwneg106_73 in106 sn73 3183.098862
Rwneg106_74 in106 sn74 11140.846016
Rwneg106_75 in106 sn75 11140.846016
Rwneg106_76 in106 sn76 11140.846016
Rwneg106_77 in106 sn77 3183.098862
Rwneg106_78 in106 sn78 3183.098862
Rwneg106_79 in106 sn79 11140.846016
Rwneg106_80 in106 sn80 3183.098862
Rwneg106_81 in106 sn81 3183.098862
Rwneg106_82 in106 sn82 11140.846016
Rwneg106_83 in106 sn83 3183.098862
Rwneg106_84 in106 sn84 11140.846016
Rwneg106_85 in106 sn85 3183.098862
Rwneg106_86 in106 sn86 11140.846016
Rwneg106_87 in106 sn87 11140.846016
Rwneg106_88 in106 sn88 11140.846016
Rwneg106_89 in106 sn89 3183.098862
Rwneg106_90 in106 sn90 3183.098862
Rwneg106_91 in106 sn91 3183.098862
Rwneg106_92 in106 sn92 11140.846016
Rwneg106_93 in106 sn93 11140.846016
Rwneg106_94 in106 sn94 3183.098862
Rwneg106_95 in106 sn95 3183.098862
Rwneg106_96 in106 sn96 11140.846016
Rwneg106_97 in106 sn97 11140.846016
Rwneg106_98 in106 sn98 11140.846016
Rwneg106_99 in106 sn99 3183.098862
Rwneg106_100 in106 sn100 3183.098862
Rwneg107_1 in107 sn1 11140.846016
Rwneg107_2 in107 sn2 3183.098862
Rwneg107_3 in107 sn3 11140.846016
Rwneg107_4 in107 sn4 11140.846016
Rwneg107_5 in107 sn5 3183.098862
Rwneg107_6 in107 sn6 11140.846016
Rwneg107_7 in107 sn7 11140.846016
Rwneg107_8 in107 sn8 11140.846016
Rwneg107_9 in107 sn9 11140.846016
Rwneg107_10 in107 sn10 3183.098862
Rwneg107_11 in107 sn11 3183.098862
Rwneg107_12 in107 sn12 11140.846016
Rwneg107_13 in107 sn13 11140.846016
Rwneg107_14 in107 sn14 11140.846016
Rwneg107_15 in107 sn15 11140.846016
Rwneg107_16 in107 sn16 11140.846016
Rwneg107_17 in107 sn17 3183.098862
Rwneg107_18 in107 sn18 11140.846016
Rwneg107_19 in107 sn19 11140.846016
Rwneg107_20 in107 sn20 3183.098862
Rwneg107_21 in107 sn21 3183.098862
Rwneg107_22 in107 sn22 3183.098862
Rwneg107_23 in107 sn23 11140.846016
Rwneg107_24 in107 sn24 11140.846016
Rwneg107_25 in107 sn25 11140.846016
Rwneg107_26 in107 sn26 3183.098862
Rwneg107_27 in107 sn27 3183.098862
Rwneg107_28 in107 sn28 11140.846016
Rwneg107_29 in107 sn29 11140.846016
Rwneg107_30 in107 sn30 11140.846016
Rwneg107_31 in107 sn31 11140.846016
Rwneg107_32 in107 sn32 3183.098862
Rwneg107_33 in107 sn33 3183.098862
Rwneg107_34 in107 sn34 3183.098862
Rwneg107_35 in107 sn35 11140.846016
Rwneg107_36 in107 sn36 11140.846016
Rwneg107_37 in107 sn37 11140.846016
Rwneg107_38 in107 sn38 11140.846016
Rwneg107_39 in107 sn39 11140.846016
Rwneg107_40 in107 sn40 11140.846016
Rwneg107_41 in107 sn41 11140.846016
Rwneg107_42 in107 sn42 3183.098862
Rwneg107_43 in107 sn43 3183.098862
Rwneg107_44 in107 sn44 3183.098862
Rwneg107_45 in107 sn45 11140.846016
Rwneg107_46 in107 sn46 11140.846016
Rwneg107_47 in107 sn47 11140.846016
Rwneg107_48 in107 sn48 3183.098862
Rwneg107_49 in107 sn49 3183.098862
Rwneg107_50 in107 sn50 3183.098862
Rwneg107_51 in107 sn51 3183.098862
Rwneg107_52 in107 sn52 3183.098862
Rwneg107_53 in107 sn53 3183.098862
Rwneg107_54 in107 sn54 3183.098862
Rwneg107_55 in107 sn55 11140.846016
Rwneg107_56 in107 sn56 3183.098862
Rwneg107_57 in107 sn57 11140.846016
Rwneg107_58 in107 sn58 3183.098862
Rwneg107_59 in107 sn59 3183.098862
Rwneg107_60 in107 sn60 11140.846016
Rwneg107_61 in107 sn61 11140.846016
Rwneg107_62 in107 sn62 11140.846016
Rwneg107_63 in107 sn63 3183.098862
Rwneg107_64 in107 sn64 3183.098862
Rwneg107_65 in107 sn65 3183.098862
Rwneg107_66 in107 sn66 3183.098862
Rwneg107_67 in107 sn67 11140.846016
Rwneg107_68 in107 sn68 3183.098862
Rwneg107_69 in107 sn69 11140.846016
Rwneg107_70 in107 sn70 3183.098862
Rwneg107_71 in107 sn71 11140.846016
Rwneg107_72 in107 sn72 3183.098862
Rwneg107_73 in107 sn73 3183.098862
Rwneg107_74 in107 sn74 11140.846016
Rwneg107_75 in107 sn75 3183.098862
Rwneg107_76 in107 sn76 11140.846016
Rwneg107_77 in107 sn77 3183.098862
Rwneg107_78 in107 sn78 11140.846016
Rwneg107_79 in107 sn79 11140.846016
Rwneg107_80 in107 sn80 11140.846016
Rwneg107_81 in107 sn81 3183.098862
Rwneg107_82 in107 sn82 3183.098862
Rwneg107_83 in107 sn83 3183.098862
Rwneg107_84 in107 sn84 3183.098862
Rwneg107_85 in107 sn85 3183.098862
Rwneg107_86 in107 sn86 3183.098862
Rwneg107_87 in107 sn87 11140.846016
Rwneg107_88 in107 sn88 11140.846016
Rwneg107_89 in107 sn89 11140.846016
Rwneg107_90 in107 sn90 3183.098862
Rwneg107_91 in107 sn91 3183.098862
Rwneg107_92 in107 sn92 3183.098862
Rwneg107_93 in107 sn93 3183.098862
Rwneg107_94 in107 sn94 3183.098862
Rwneg107_95 in107 sn95 11140.846016
Rwneg107_96 in107 sn96 3183.098862
Rwneg107_97 in107 sn97 3183.098862
Rwneg107_98 in107 sn98 3183.098862
Rwneg107_99 in107 sn99 11140.846016
Rwneg107_100 in107 sn100 3183.098862
Rwneg108_1 in108 sn1 11140.846016
Rwneg108_2 in108 sn2 11140.846016
Rwneg108_3 in108 sn3 3183.098862
Rwneg108_4 in108 sn4 3183.098862
Rwneg108_5 in108 sn5 11140.846016
Rwneg108_6 in108 sn6 11140.846016
Rwneg108_7 in108 sn7 11140.846016
Rwneg108_8 in108 sn8 11140.846016
Rwneg108_9 in108 sn9 11140.846016
Rwneg108_10 in108 sn10 11140.846016
Rwneg108_11 in108 sn11 3183.098862
Rwneg108_12 in108 sn12 11140.846016
Rwneg108_13 in108 sn13 3183.098862
Rwneg108_14 in108 sn14 3183.098862
Rwneg108_15 in108 sn15 11140.846016
Rwneg108_16 in108 sn16 11140.846016
Rwneg108_17 in108 sn17 3183.098862
Rwneg108_18 in108 sn18 3183.098862
Rwneg108_19 in108 sn19 3183.098862
Rwneg108_20 in108 sn20 3183.098862
Rwneg108_21 in108 sn21 11140.846016
Rwneg108_22 in108 sn22 11140.846016
Rwneg108_23 in108 sn23 11140.846016
Rwneg108_24 in108 sn24 3183.098862
Rwneg108_25 in108 sn25 11140.846016
Rwneg108_26 in108 sn26 11140.846016
Rwneg108_27 in108 sn27 11140.846016
Rwneg108_28 in108 sn28 3183.098862
Rwneg108_29 in108 sn29 11140.846016
Rwneg108_30 in108 sn30 11140.846016
Rwneg108_31 in108 sn31 11140.846016
Rwneg108_32 in108 sn32 3183.098862
Rwneg108_33 in108 sn33 11140.846016
Rwneg108_34 in108 sn34 3183.098862
Rwneg108_35 in108 sn35 11140.846016
Rwneg108_36 in108 sn36 11140.846016
Rwneg108_37 in108 sn37 11140.846016
Rwneg108_38 in108 sn38 11140.846016
Rwneg108_39 in108 sn39 11140.846016
Rwneg108_40 in108 sn40 3183.098862
Rwneg108_41 in108 sn41 3183.098862
Rwneg108_42 in108 sn42 11140.846016
Rwneg108_43 in108 sn43 3183.098862
Rwneg108_44 in108 sn44 11140.846016
Rwneg108_45 in108 sn45 11140.846016
Rwneg108_46 in108 sn46 3183.098862
Rwneg108_47 in108 sn47 3183.098862
Rwneg108_48 in108 sn48 11140.846016
Rwneg108_49 in108 sn49 11140.846016
Rwneg108_50 in108 sn50 11140.846016
Rwneg108_51 in108 sn51 11140.846016
Rwneg108_52 in108 sn52 3183.098862
Rwneg108_53 in108 sn53 11140.846016
Rwneg108_54 in108 sn54 3183.098862
Rwneg108_55 in108 sn55 3183.098862
Rwneg108_56 in108 sn56 11140.846016
Rwneg108_57 in108 sn57 11140.846016
Rwneg108_58 in108 sn58 11140.846016
Rwneg108_59 in108 sn59 3183.098862
Rwneg108_60 in108 sn60 3183.098862
Rwneg108_61 in108 sn61 11140.846016
Rwneg108_62 in108 sn62 3183.098862
Rwneg108_63 in108 sn63 3183.098862
Rwneg108_64 in108 sn64 11140.846016
Rwneg108_65 in108 sn65 3183.098862
Rwneg108_66 in108 sn66 3183.098862
Rwneg108_67 in108 sn67 11140.846016
Rwneg108_68 in108 sn68 3183.098862
Rwneg108_69 in108 sn69 11140.846016
Rwneg108_70 in108 sn70 3183.098862
Rwneg108_71 in108 sn71 11140.846016
Rwneg108_72 in108 sn72 11140.846016
Rwneg108_73 in108 sn73 11140.846016
Rwneg108_74 in108 sn74 3183.098862
Rwneg108_75 in108 sn75 3183.098862
Rwneg108_76 in108 sn76 11140.846016
Rwneg108_77 in108 sn77 11140.846016
Rwneg108_78 in108 sn78 3183.098862
Rwneg108_79 in108 sn79 11140.846016
Rwneg108_80 in108 sn80 3183.098862
Rwneg108_81 in108 sn81 11140.846016
Rwneg108_82 in108 sn82 3183.098862
Rwneg108_83 in108 sn83 3183.098862
Rwneg108_84 in108 sn84 3183.098862
Rwneg108_85 in108 sn85 11140.846016
Rwneg108_86 in108 sn86 11140.846016
Rwneg108_87 in108 sn87 3183.098862
Rwneg108_88 in108 sn88 11140.846016
Rwneg108_89 in108 sn89 3183.098862
Rwneg108_90 in108 sn90 3183.098862
Rwneg108_91 in108 sn91 11140.846016
Rwneg108_92 in108 sn92 3183.098862
Rwneg108_93 in108 sn93 3183.098862
Rwneg108_94 in108 sn94 11140.846016
Rwneg108_95 in108 sn95 3183.098862
Rwneg108_96 in108 sn96 3183.098862
Rwneg108_97 in108 sn97 11140.846016
Rwneg108_98 in108 sn98 3183.098862
Rwneg108_99 in108 sn99 11140.846016
Rwneg108_100 in108 sn100 3183.098862
Rwneg109_1 in109 sn1 3183.098862
Rwneg109_2 in109 sn2 3183.098862
Rwneg109_3 in109 sn3 3183.098862
Rwneg109_4 in109 sn4 3183.098862
Rwneg109_5 in109 sn5 11140.846016
Rwneg109_6 in109 sn6 11140.846016
Rwneg109_7 in109 sn7 11140.846016
Rwneg109_8 in109 sn8 11140.846016
Rwneg109_9 in109 sn9 3183.098862
Rwneg109_10 in109 sn10 11140.846016
Rwneg109_11 in109 sn11 11140.846016
Rwneg109_12 in109 sn12 11140.846016
Rwneg109_13 in109 sn13 3183.098862
Rwneg109_14 in109 sn14 3183.098862
Rwneg109_15 in109 sn15 11140.846016
Rwneg109_16 in109 sn16 11140.846016
Rwneg109_17 in109 sn17 3183.098862
Rwneg109_18 in109 sn18 3183.098862
Rwneg109_19 in109 sn19 3183.098862
Rwneg109_20 in109 sn20 3183.098862
Rwneg109_21 in109 sn21 11140.846016
Rwneg109_22 in109 sn22 3183.098862
Rwneg109_23 in109 sn23 3183.098862
Rwneg109_24 in109 sn24 3183.098862
Rwneg109_25 in109 sn25 11140.846016
Rwneg109_26 in109 sn26 11140.846016
Rwneg109_27 in109 sn27 11140.846016
Rwneg109_28 in109 sn28 3183.098862
Rwneg109_29 in109 sn29 3183.098862
Rwneg109_30 in109 sn30 3183.098862
Rwneg109_31 in109 sn31 11140.846016
Rwneg109_32 in109 sn32 11140.846016
Rwneg109_33 in109 sn33 3183.098862
Rwneg109_34 in109 sn34 11140.846016
Rwneg109_35 in109 sn35 11140.846016
Rwneg109_36 in109 sn36 3183.098862
Rwneg109_37 in109 sn37 3183.098862
Rwneg109_38 in109 sn38 11140.846016
Rwneg109_39 in109 sn39 11140.846016
Rwneg109_40 in109 sn40 11140.846016
Rwneg109_41 in109 sn41 3183.098862
Rwneg109_42 in109 sn42 3183.098862
Rwneg109_43 in109 sn43 3183.098862
Rwneg109_44 in109 sn44 11140.846016
Rwneg109_45 in109 sn45 11140.846016
Rwneg109_46 in109 sn46 11140.846016
Rwneg109_47 in109 sn47 3183.098862
Rwneg109_48 in109 sn48 3183.098862
Rwneg109_49 in109 sn49 3183.098862
Rwneg109_50 in109 sn50 3183.098862
Rwneg109_51 in109 sn51 3183.098862
Rwneg109_52 in109 sn52 3183.098862
Rwneg109_53 in109 sn53 11140.846016
Rwneg109_54 in109 sn54 3183.098862
Rwneg109_55 in109 sn55 3183.098862
Rwneg109_56 in109 sn56 11140.846016
Rwneg109_57 in109 sn57 11140.846016
Rwneg109_58 in109 sn58 3183.098862
Rwneg109_59 in109 sn59 3183.098862
Rwneg109_60 in109 sn60 11140.846016
Rwneg109_61 in109 sn61 11140.846016
Rwneg109_62 in109 sn62 11140.846016
Rwneg109_63 in109 sn63 3183.098862
Rwneg109_64 in109 sn64 3183.098862
Rwneg109_65 in109 sn65 3183.098862
Rwneg109_66 in109 sn66 11140.846016
Rwneg109_67 in109 sn67 3183.098862
Rwneg109_68 in109 sn68 11140.846016
Rwneg109_69 in109 sn69 3183.098862
Rwneg109_70 in109 sn70 3183.098862
Rwneg109_71 in109 sn71 11140.846016
Rwneg109_72 in109 sn72 11140.846016
Rwneg109_73 in109 sn73 3183.098862
Rwneg109_74 in109 sn74 3183.098862
Rwneg109_75 in109 sn75 3183.098862
Rwneg109_76 in109 sn76 11140.846016
Rwneg109_77 in109 sn77 11140.846016
Rwneg109_78 in109 sn78 11140.846016
Rwneg109_79 in109 sn79 11140.846016
Rwneg109_80 in109 sn80 11140.846016
Rwneg109_81 in109 sn81 3183.098862
Rwneg109_82 in109 sn82 11140.846016
Rwneg109_83 in109 sn83 11140.846016
Rwneg109_84 in109 sn84 3183.098862
Rwneg109_85 in109 sn85 11140.846016
Rwneg109_86 in109 sn86 3183.098862
Rwneg109_87 in109 sn87 11140.846016
Rwneg109_88 in109 sn88 3183.098862
Rwneg109_89 in109 sn89 11140.846016
Rwneg109_90 in109 sn90 3183.098862
Rwneg109_91 in109 sn91 3183.098862
Rwneg109_92 in109 sn92 11140.846016
Rwneg109_93 in109 sn93 11140.846016
Rwneg109_94 in109 sn94 11140.846016
Rwneg109_95 in109 sn95 3183.098862
Rwneg109_96 in109 sn96 3183.098862
Rwneg109_97 in109 sn97 3183.098862
Rwneg109_98 in109 sn98 3183.098862
Rwneg109_99 in109 sn99 3183.098862
Rwneg109_100 in109 sn100 11140.846016
Rwneg110_1 in110 sn1 3183.098862
Rwneg110_2 in110 sn2 3183.098862
Rwneg110_3 in110 sn3 3183.098862
Rwneg110_4 in110 sn4 3183.098862
Rwneg110_5 in110 sn5 3183.098862
Rwneg110_6 in110 sn6 11140.846016
Rwneg110_7 in110 sn7 11140.846016
Rwneg110_8 in110 sn8 11140.846016
Rwneg110_9 in110 sn9 3183.098862
Rwneg110_10 in110 sn10 11140.846016
Rwneg110_11 in110 sn11 3183.098862
Rwneg110_12 in110 sn12 11140.846016
Rwneg110_13 in110 sn13 3183.098862
Rwneg110_14 in110 sn14 11140.846016
Rwneg110_15 in110 sn15 11140.846016
Rwneg110_16 in110 sn16 3183.098862
Rwneg110_17 in110 sn17 3183.098862
Rwneg110_18 in110 sn18 3183.098862
Rwneg110_19 in110 sn19 11140.846016
Rwneg110_20 in110 sn20 11140.846016
Rwneg110_21 in110 sn21 3183.098862
Rwneg110_22 in110 sn22 11140.846016
Rwneg110_23 in110 sn23 11140.846016
Rwneg110_24 in110 sn24 11140.846016
Rwneg110_25 in110 sn25 11140.846016
Rwneg110_26 in110 sn26 11140.846016
Rwneg110_27 in110 sn27 11140.846016
Rwneg110_28 in110 sn28 11140.846016
Rwneg110_29 in110 sn29 3183.098862
Rwneg110_30 in110 sn30 11140.846016
Rwneg110_31 in110 sn31 11140.846016
Rwneg110_32 in110 sn32 11140.846016
Rwneg110_33 in110 sn33 11140.846016
Rwneg110_34 in110 sn34 3183.098862
Rwneg110_35 in110 sn35 11140.846016
Rwneg110_36 in110 sn36 11140.846016
Rwneg110_37 in110 sn37 11140.846016
Rwneg110_38 in110 sn38 11140.846016
Rwneg110_39 in110 sn39 11140.846016
Rwneg110_40 in110 sn40 3183.098862
Rwneg110_41 in110 sn41 3183.098862
Rwneg110_42 in110 sn42 11140.846016
Rwneg110_43 in110 sn43 11140.846016
Rwneg110_44 in110 sn44 11140.846016
Rwneg110_45 in110 sn45 11140.846016
Rwneg110_46 in110 sn46 11140.846016
Rwneg110_47 in110 sn47 11140.846016
Rwneg110_48 in110 sn48 11140.846016
Rwneg110_49 in110 sn49 3183.098862
Rwneg110_50 in110 sn50 3183.098862
Rwneg110_51 in110 sn51 3183.098862
Rwneg110_52 in110 sn52 11140.846016
Rwneg110_53 in110 sn53 11140.846016
Rwneg110_54 in110 sn54 11140.846016
Rwneg110_55 in110 sn55 11140.846016
Rwneg110_56 in110 sn56 11140.846016
Rwneg110_57 in110 sn57 11140.846016
Rwneg110_58 in110 sn58 3183.098862
Rwneg110_59 in110 sn59 3183.098862
Rwneg110_60 in110 sn60 11140.846016
Rwneg110_61 in110 sn61 3183.098862
Rwneg110_62 in110 sn62 11140.846016
Rwneg110_63 in110 sn63 3183.098862
Rwneg110_64 in110 sn64 11140.846016
Rwneg110_65 in110 sn65 11140.846016
Rwneg110_66 in110 sn66 3183.098862
Rwneg110_67 in110 sn67 11140.846016
Rwneg110_68 in110 sn68 11140.846016
Rwneg110_69 in110 sn69 11140.846016
Rwneg110_70 in110 sn70 11140.846016
Rwneg110_71 in110 sn71 3183.098862
Rwneg110_72 in110 sn72 3183.098862
Rwneg110_73 in110 sn73 3183.098862
Rwneg110_74 in110 sn74 11140.846016
Rwneg110_75 in110 sn75 11140.846016
Rwneg110_76 in110 sn76 11140.846016
Rwneg110_77 in110 sn77 3183.098862
Rwneg110_78 in110 sn78 11140.846016
Rwneg110_79 in110 sn79 11140.846016
Rwneg110_80 in110 sn80 3183.098862
Rwneg110_81 in110 sn81 3183.098862
Rwneg110_82 in110 sn82 11140.846016
Rwneg110_83 in110 sn83 11140.846016
Rwneg110_84 in110 sn84 11140.846016
Rwneg110_85 in110 sn85 3183.098862
Rwneg110_86 in110 sn86 11140.846016
Rwneg110_87 in110 sn87 11140.846016
Rwneg110_88 in110 sn88 11140.846016
Rwneg110_89 in110 sn89 3183.098862
Rwneg110_90 in110 sn90 3183.098862
Rwneg110_91 in110 sn91 11140.846016
Rwneg110_92 in110 sn92 11140.846016
Rwneg110_93 in110 sn93 3183.098862
Rwneg110_94 in110 sn94 11140.846016
Rwneg110_95 in110 sn95 3183.098862
Rwneg110_96 in110 sn96 11140.846016
Rwneg110_97 in110 sn97 3183.098862
Rwneg110_98 in110 sn98 11140.846016
Rwneg110_99 in110 sn99 11140.846016
Rwneg110_100 in110 sn100 3183.098862
Rwneg111_1 in111 sn1 11140.846016
Rwneg111_2 in111 sn2 11140.846016
Rwneg111_3 in111 sn3 11140.846016
Rwneg111_4 in111 sn4 11140.846016
Rwneg111_5 in111 sn5 3183.098862
Rwneg111_6 in111 sn6 11140.846016
Rwneg111_7 in111 sn7 11140.846016
Rwneg111_8 in111 sn8 11140.846016
Rwneg111_9 in111 sn9 3183.098862
Rwneg111_10 in111 sn10 11140.846016
Rwneg111_11 in111 sn11 3183.098862
Rwneg111_12 in111 sn12 11140.846016
Rwneg111_13 in111 sn13 11140.846016
Rwneg111_14 in111 sn14 11140.846016
Rwneg111_15 in111 sn15 11140.846016
Rwneg111_16 in111 sn16 11140.846016
Rwneg111_17 in111 sn17 11140.846016
Rwneg111_18 in111 sn18 11140.846016
Rwneg111_19 in111 sn19 11140.846016
Rwneg111_20 in111 sn20 11140.846016
Rwneg111_21 in111 sn21 3183.098862
Rwneg111_22 in111 sn22 3183.098862
Rwneg111_23 in111 sn23 3183.098862
Rwneg111_24 in111 sn24 11140.846016
Rwneg111_25 in111 sn25 11140.846016
Rwneg111_26 in111 sn26 11140.846016
Rwneg111_27 in111 sn27 3183.098862
Rwneg111_28 in111 sn28 3183.098862
Rwneg111_29 in111 sn29 3183.098862
Rwneg111_30 in111 sn30 11140.846016
Rwneg111_31 in111 sn31 11140.846016
Rwneg111_32 in111 sn32 11140.846016
Rwneg111_33 in111 sn33 11140.846016
Rwneg111_34 in111 sn34 11140.846016
Rwneg111_35 in111 sn35 3183.098862
Rwneg111_36 in111 sn36 3183.098862
Rwneg111_37 in111 sn37 3183.098862
Rwneg111_38 in111 sn38 3183.098862
Rwneg111_39 in111 sn39 11140.846016
Rwneg111_40 in111 sn40 11140.846016
Rwneg111_41 in111 sn41 11140.846016
Rwneg111_42 in111 sn42 11140.846016
Rwneg111_43 in111 sn43 3183.098862
Rwneg111_44 in111 sn44 11140.846016
Rwneg111_45 in111 sn45 3183.098862
Rwneg111_46 in111 sn46 11140.846016
Rwneg111_47 in111 sn47 3183.098862
Rwneg111_48 in111 sn48 3183.098862
Rwneg111_49 in111 sn49 11140.846016
Rwneg111_50 in111 sn50 11140.846016
Rwneg111_51 in111 sn51 11140.846016
Rwneg111_52 in111 sn52 11140.846016
Rwneg111_53 in111 sn53 11140.846016
Rwneg111_54 in111 sn54 3183.098862
Rwneg111_55 in111 sn55 3183.098862
Rwneg111_56 in111 sn56 11140.846016
Rwneg111_57 in111 sn57 11140.846016
Rwneg111_58 in111 sn58 11140.846016
Rwneg111_59 in111 sn59 3183.098862
Rwneg111_60 in111 sn60 11140.846016
Rwneg111_61 in111 sn61 3183.098862
Rwneg111_62 in111 sn62 11140.846016
Rwneg111_63 in111 sn63 3183.098862
Rwneg111_64 in111 sn64 3183.098862
Rwneg111_65 in111 sn65 11140.846016
Rwneg111_66 in111 sn66 11140.846016
Rwneg111_67 in111 sn67 11140.846016
Rwneg111_68 in111 sn68 11140.846016
Rwneg111_69 in111 sn69 11140.846016
Rwneg111_70 in111 sn70 11140.846016
Rwneg111_71 in111 sn71 3183.098862
Rwneg111_72 in111 sn72 11140.846016
Rwneg111_73 in111 sn73 3183.098862
Rwneg111_74 in111 sn74 11140.846016
Rwneg111_75 in111 sn75 3183.098862
Rwneg111_76 in111 sn76 11140.846016
Rwneg111_77 in111 sn77 3183.098862
Rwneg111_78 in111 sn78 11140.846016
Rwneg111_79 in111 sn79 3183.098862
Rwneg111_80 in111 sn80 3183.098862
Rwneg111_81 in111 sn81 3183.098862
Rwneg111_82 in111 sn82 3183.098862
Rwneg111_83 in111 sn83 11140.846016
Rwneg111_84 in111 sn84 3183.098862
Rwneg111_85 in111 sn85 3183.098862
Rwneg111_86 in111 sn86 3183.098862
Rwneg111_87 in111 sn87 3183.098862
Rwneg111_88 in111 sn88 11140.846016
Rwneg111_89 in111 sn89 11140.846016
Rwneg111_90 in111 sn90 3183.098862
Rwneg111_91 in111 sn91 3183.098862
Rwneg111_92 in111 sn92 11140.846016
Rwneg111_93 in111 sn93 3183.098862
Rwneg111_94 in111 sn94 11140.846016
Rwneg111_95 in111 sn95 3183.098862
Rwneg111_96 in111 sn96 3183.098862
Rwneg111_97 in111 sn97 3183.098862
Rwneg111_98 in111 sn98 11140.846016
Rwneg111_99 in111 sn99 11140.846016
Rwneg111_100 in111 sn100 11140.846016
Rwneg112_1 in112 sn1 11140.846016
Rwneg112_2 in112 sn2 11140.846016
Rwneg112_3 in112 sn3 3183.098862
Rwneg112_4 in112 sn4 3183.098862
Rwneg112_5 in112 sn5 3183.098862
Rwneg112_6 in112 sn6 11140.846016
Rwneg112_7 in112 sn7 3183.098862
Rwneg112_8 in112 sn8 3183.098862
Rwneg112_9 in112 sn9 11140.846016
Rwneg112_10 in112 sn10 11140.846016
Rwneg112_11 in112 sn11 3183.098862
Rwneg112_12 in112 sn12 11140.846016
Rwneg112_13 in112 sn13 3183.098862
Rwneg112_14 in112 sn14 11140.846016
Rwneg112_15 in112 sn15 11140.846016
Rwneg112_16 in112 sn16 3183.098862
Rwneg112_17 in112 sn17 3183.098862
Rwneg112_18 in112 sn18 3183.098862
Rwneg112_19 in112 sn19 11140.846016
Rwneg112_20 in112 sn20 11140.846016
Rwneg112_21 in112 sn21 3183.098862
Rwneg112_22 in112 sn22 11140.846016
Rwneg112_23 in112 sn23 3183.098862
Rwneg112_24 in112 sn24 11140.846016
Rwneg112_25 in112 sn25 11140.846016
Rwneg112_26 in112 sn26 11140.846016
Rwneg112_27 in112 sn27 11140.846016
Rwneg112_28 in112 sn28 3183.098862
Rwneg112_29 in112 sn29 3183.098862
Rwneg112_30 in112 sn30 11140.846016
Rwneg112_31 in112 sn31 11140.846016
Rwneg112_32 in112 sn32 11140.846016
Rwneg112_33 in112 sn33 3183.098862
Rwneg112_34 in112 sn34 11140.846016
Rwneg112_35 in112 sn35 11140.846016
Rwneg112_36 in112 sn36 3183.098862
Rwneg112_37 in112 sn37 3183.098862
Rwneg112_38 in112 sn38 3183.098862
Rwneg112_39 in112 sn39 3183.098862
Rwneg112_40 in112 sn40 3183.098862
Rwneg112_41 in112 sn41 11140.846016
Rwneg112_42 in112 sn42 3183.098862
Rwneg112_43 in112 sn43 11140.846016
Rwneg112_44 in112 sn44 11140.846016
Rwneg112_45 in112 sn45 3183.098862
Rwneg112_46 in112 sn46 3183.098862
Rwneg112_47 in112 sn47 3183.098862
Rwneg112_48 in112 sn48 3183.098862
Rwneg112_49 in112 sn49 11140.846016
Rwneg112_50 in112 sn50 3183.098862
Rwneg112_51 in112 sn51 11140.846016
Rwneg112_52 in112 sn52 3183.098862
Rwneg112_53 in112 sn53 3183.098862
Rwneg112_54 in112 sn54 3183.098862
Rwneg112_55 in112 sn55 3183.098862
Rwneg112_56 in112 sn56 11140.846016
Rwneg112_57 in112 sn57 11140.846016
Rwneg112_58 in112 sn58 11140.846016
Rwneg112_59 in112 sn59 3183.098862
Rwneg112_60 in112 sn60 3183.098862
Rwneg112_61 in112 sn61 3183.098862
Rwneg112_62 in112 sn62 11140.846016
Rwneg112_63 in112 sn63 11140.846016
Rwneg112_64 in112 sn64 11140.846016
Rwneg112_65 in112 sn65 11140.846016
Rwneg112_66 in112 sn66 3183.098862
Rwneg112_67 in112 sn67 11140.846016
Rwneg112_68 in112 sn68 3183.098862
Rwneg112_69 in112 sn69 3183.098862
Rwneg112_70 in112 sn70 3183.098862
Rwneg112_71 in112 sn71 3183.098862
Rwneg112_72 in112 sn72 11140.846016
Rwneg112_73 in112 sn73 3183.098862
Rwneg112_74 in112 sn74 3183.098862
Rwneg112_75 in112 sn75 3183.098862
Rwneg112_76 in112 sn76 3183.098862
Rwneg112_77 in112 sn77 3183.098862
Rwneg112_78 in112 sn78 3183.098862
Rwneg112_79 in112 sn79 3183.098862
Rwneg112_80 in112 sn80 11140.846016
Rwneg112_81 in112 sn81 11140.846016
Rwneg112_82 in112 sn82 11140.846016
Rwneg112_83 in112 sn83 11140.846016
Rwneg112_84 in112 sn84 11140.846016
Rwneg112_85 in112 sn85 11140.846016
Rwneg112_86 in112 sn86 11140.846016
Rwneg112_87 in112 sn87 3183.098862
Rwneg112_88 in112 sn88 3183.098862
Rwneg112_89 in112 sn89 11140.846016
Rwneg112_90 in112 sn90 3183.098862
Rwneg112_91 in112 sn91 11140.846016
Rwneg112_92 in112 sn92 11140.846016
Rwneg112_93 in112 sn93 11140.846016
Rwneg112_94 in112 sn94 3183.098862
Rwneg112_95 in112 sn95 3183.098862
Rwneg112_96 in112 sn96 3183.098862
Rwneg112_97 in112 sn97 11140.846016
Rwneg112_98 in112 sn98 11140.846016
Rwneg112_99 in112 sn99 11140.846016
Rwneg112_100 in112 sn100 11140.846016
Rwneg113_1 in113 sn1 11140.846016
Rwneg113_2 in113 sn2 11140.846016
Rwneg113_3 in113 sn3 3183.098862
Rwneg113_4 in113 sn4 3183.098862
Rwneg113_5 in113 sn5 3183.098862
Rwneg113_6 in113 sn6 3183.098862
Rwneg113_7 in113 sn7 11140.846016
Rwneg113_8 in113 sn8 11140.846016
Rwneg113_9 in113 sn9 11140.846016
Rwneg113_10 in113 sn10 11140.846016
Rwneg113_11 in113 sn11 11140.846016
Rwneg113_12 in113 sn12 3183.098862
Rwneg113_13 in113 sn13 11140.846016
Rwneg113_14 in113 sn14 3183.098862
Rwneg113_15 in113 sn15 3183.098862
Rwneg113_16 in113 sn16 3183.098862
Rwneg113_17 in113 sn17 3183.098862
Rwneg113_18 in113 sn18 11140.846016
Rwneg113_19 in113 sn19 3183.098862
Rwneg113_20 in113 sn20 11140.846016
Rwneg113_21 in113 sn21 11140.846016
Rwneg113_22 in113 sn22 3183.098862
Rwneg113_23 in113 sn23 3183.098862
Rwneg113_24 in113 sn24 11140.846016
Rwneg113_25 in113 sn25 3183.098862
Rwneg113_26 in113 sn26 3183.098862
Rwneg113_27 in113 sn27 11140.846016
Rwneg113_28 in113 sn28 3183.098862
Rwneg113_29 in113 sn29 11140.846016
Rwneg113_30 in113 sn30 3183.098862
Rwneg113_31 in113 sn31 3183.098862
Rwneg113_32 in113 sn32 3183.098862
Rwneg113_33 in113 sn33 3183.098862
Rwneg113_34 in113 sn34 11140.846016
Rwneg113_35 in113 sn35 11140.846016
Rwneg113_36 in113 sn36 3183.098862
Rwneg113_37 in113 sn37 3183.098862
Rwneg113_38 in113 sn38 3183.098862
Rwneg113_39 in113 sn39 3183.098862
Rwneg113_40 in113 sn40 3183.098862
Rwneg113_41 in113 sn41 11140.846016
Rwneg113_42 in113 sn42 11140.846016
Rwneg113_43 in113 sn43 11140.846016
Rwneg113_44 in113 sn44 3183.098862
Rwneg113_45 in113 sn45 3183.098862
Rwneg113_46 in113 sn46 3183.098862
Rwneg113_47 in113 sn47 3183.098862
Rwneg113_48 in113 sn48 3183.098862
Rwneg113_49 in113 sn49 3183.098862
Rwneg113_50 in113 sn50 3183.098862
Rwneg113_51 in113 sn51 3183.098862
Rwneg113_52 in113 sn52 11140.846016
Rwneg113_53 in113 sn53 11140.846016
Rwneg113_54 in113 sn54 11140.846016
Rwneg113_55 in113 sn55 3183.098862
Rwneg113_56 in113 sn56 3183.098862
Rwneg113_57 in113 sn57 3183.098862
Rwneg113_58 in113 sn58 3183.098862
Rwneg113_59 in113 sn59 11140.846016
Rwneg113_60 in113 sn60 11140.846016
Rwneg113_61 in113 sn61 3183.098862
Rwneg113_62 in113 sn62 11140.846016
Rwneg113_63 in113 sn63 3183.098862
Rwneg113_64 in113 sn64 11140.846016
Rwneg113_65 in113 sn65 11140.846016
Rwneg113_66 in113 sn66 3183.098862
Rwneg113_67 in113 sn67 3183.098862
Rwneg113_68 in113 sn68 3183.098862
Rwneg113_69 in113 sn69 3183.098862
Rwneg113_70 in113 sn70 11140.846016
Rwneg113_71 in113 sn71 11140.846016
Rwneg113_72 in113 sn72 3183.098862
Rwneg113_73 in113 sn73 3183.098862
Rwneg113_74 in113 sn74 11140.846016
Rwneg113_75 in113 sn75 3183.098862
Rwneg113_76 in113 sn76 11140.846016
Rwneg113_77 in113 sn77 3183.098862
Rwneg113_78 in113 sn78 11140.846016
Rwneg113_79 in113 sn79 3183.098862
Rwneg113_80 in113 sn80 3183.098862
Rwneg113_81 in113 sn81 3183.098862
Rwneg113_82 in113 sn82 3183.098862
Rwneg113_83 in113 sn83 3183.098862
Rwneg113_84 in113 sn84 3183.098862
Rwneg113_85 in113 sn85 3183.098862
Rwneg113_86 in113 sn86 11140.846016
Rwneg113_87 in113 sn87 11140.846016
Rwneg113_88 in113 sn88 11140.846016
Rwneg113_89 in113 sn89 3183.098862
Rwneg113_90 in113 sn90 11140.846016
Rwneg113_91 in113 sn91 11140.846016
Rwneg113_92 in113 sn92 11140.846016
Rwneg113_93 in113 sn93 11140.846016
Rwneg113_94 in113 sn94 3183.098862
Rwneg113_95 in113 sn95 3183.098862
Rwneg113_96 in113 sn96 3183.098862
Rwneg113_97 in113 sn97 3183.098862
Rwneg113_98 in113 sn98 11140.846016
Rwneg113_99 in113 sn99 3183.098862
Rwneg113_100 in113 sn100 11140.846016
Rwneg114_1 in114 sn1 11140.846016
Rwneg114_2 in114 sn2 11140.846016
Rwneg114_3 in114 sn3 3183.098862
Rwneg114_4 in114 sn4 11140.846016
Rwneg114_5 in114 sn5 3183.098862
Rwneg114_6 in114 sn6 11140.846016
Rwneg114_7 in114 sn7 11140.846016
Rwneg114_8 in114 sn8 11140.846016
Rwneg114_9 in114 sn9 11140.846016
Rwneg114_10 in114 sn10 3183.098862
Rwneg114_11 in114 sn11 3183.098862
Rwneg114_12 in114 sn12 11140.846016
Rwneg114_13 in114 sn13 3183.098862
Rwneg114_14 in114 sn14 11140.846016
Rwneg114_15 in114 sn15 3183.098862
Rwneg114_16 in114 sn16 11140.846016
Rwneg114_17 in114 sn17 11140.846016
Rwneg114_18 in114 sn18 3183.098862
Rwneg114_19 in114 sn19 11140.846016
Rwneg114_20 in114 sn20 11140.846016
Rwneg114_21 in114 sn21 3183.098862
Rwneg114_22 in114 sn22 11140.846016
Rwneg114_23 in114 sn23 3183.098862
Rwneg114_24 in114 sn24 3183.098862
Rwneg114_25 in114 sn25 11140.846016
Rwneg114_26 in114 sn26 11140.846016
Rwneg114_27 in114 sn27 11140.846016
Rwneg114_28 in114 sn28 11140.846016
Rwneg114_29 in114 sn29 3183.098862
Rwneg114_30 in114 sn30 11140.846016
Rwneg114_31 in114 sn31 3183.098862
Rwneg114_32 in114 sn32 3183.098862
Rwneg114_33 in114 sn33 3183.098862
Rwneg114_34 in114 sn34 3183.098862
Rwneg114_35 in114 sn35 11140.846016
Rwneg114_36 in114 sn36 3183.098862
Rwneg114_37 in114 sn37 11140.846016
Rwneg114_38 in114 sn38 11140.846016
Rwneg114_39 in114 sn39 11140.846016
Rwneg114_40 in114 sn40 11140.846016
Rwneg114_41 in114 sn41 11140.846016
Rwneg114_42 in114 sn42 11140.846016
Rwneg114_43 in114 sn43 3183.098862
Rwneg114_44 in114 sn44 11140.846016
Rwneg114_45 in114 sn45 3183.098862
Rwneg114_46 in114 sn46 11140.846016
Rwneg114_47 in114 sn47 3183.098862
Rwneg114_48 in114 sn48 3183.098862
Rwneg114_49 in114 sn49 3183.098862
Rwneg114_50 in114 sn50 11140.846016
Rwneg114_51 in114 sn51 11140.846016
Rwneg114_52 in114 sn52 3183.098862
Rwneg114_53 in114 sn53 11140.846016
Rwneg114_54 in114 sn54 11140.846016
Rwneg114_55 in114 sn55 3183.098862
Rwneg114_56 in114 sn56 11140.846016
Rwneg114_57 in114 sn57 11140.846016
Rwneg114_58 in114 sn58 11140.846016
Rwneg114_59 in114 sn59 3183.098862
Rwneg114_60 in114 sn60 11140.846016
Rwneg114_61 in114 sn61 3183.098862
Rwneg114_62 in114 sn62 11140.846016
Rwneg114_63 in114 sn63 3183.098862
Rwneg114_64 in114 sn64 3183.098862
Rwneg114_65 in114 sn65 3183.098862
Rwneg114_66 in114 sn66 3183.098862
Rwneg114_67 in114 sn67 11140.846016
Rwneg114_68 in114 sn68 3183.098862
Rwneg114_69 in114 sn69 11140.846016
Rwneg114_70 in114 sn70 11140.846016
Rwneg114_71 in114 sn71 11140.846016
Rwneg114_72 in114 sn72 11140.846016
Rwneg114_73 in114 sn73 11140.846016
Rwneg114_74 in114 sn74 11140.846016
Rwneg114_75 in114 sn75 3183.098862
Rwneg114_76 in114 sn76 11140.846016
Rwneg114_77 in114 sn77 3183.098862
Rwneg114_78 in114 sn78 11140.846016
Rwneg114_79 in114 sn79 3183.098862
Rwneg114_80 in114 sn80 3183.098862
Rwneg114_81 in114 sn81 3183.098862
Rwneg114_82 in114 sn82 11140.846016
Rwneg114_83 in114 sn83 11140.846016
Rwneg114_84 in114 sn84 11140.846016
Rwneg114_85 in114 sn85 3183.098862
Rwneg114_86 in114 sn86 11140.846016
Rwneg114_87 in114 sn87 3183.098862
Rwneg114_88 in114 sn88 11140.846016
Rwneg114_89 in114 sn89 11140.846016
Rwneg114_90 in114 sn90 11140.846016
Rwneg114_91 in114 sn91 3183.098862
Rwneg114_92 in114 sn92 11140.846016
Rwneg114_93 in114 sn93 3183.098862
Rwneg114_94 in114 sn94 11140.846016
Rwneg114_95 in114 sn95 3183.098862
Rwneg114_96 in114 sn96 3183.098862
Rwneg114_97 in114 sn97 3183.098862
Rwneg114_98 in114 sn98 11140.846016
Rwneg114_99 in114 sn99 11140.846016
Rwneg114_100 in114 sn100 3183.098862
Rwneg115_1 in115 sn1 11140.846016
Rwneg115_2 in115 sn2 11140.846016
Rwneg115_3 in115 sn3 3183.098862
Rwneg115_4 in115 sn4 11140.846016
Rwneg115_5 in115 sn5 11140.846016
Rwneg115_6 in115 sn6 11140.846016
Rwneg115_7 in115 sn7 3183.098862
Rwneg115_8 in115 sn8 3183.098862
Rwneg115_9 in115 sn9 3183.098862
Rwneg115_10 in115 sn10 11140.846016
Rwneg115_11 in115 sn11 3183.098862
Rwneg115_12 in115 sn12 3183.098862
Rwneg115_13 in115 sn13 3183.098862
Rwneg115_14 in115 sn14 11140.846016
Rwneg115_15 in115 sn15 11140.846016
Rwneg115_16 in115 sn16 3183.098862
Rwneg115_17 in115 sn17 11140.846016
Rwneg115_18 in115 sn18 11140.846016
Rwneg115_19 in115 sn19 3183.098862
Rwneg115_20 in115 sn20 11140.846016
Rwneg115_21 in115 sn21 11140.846016
Rwneg115_22 in115 sn22 11140.846016
Rwneg115_23 in115 sn23 3183.098862
Rwneg115_24 in115 sn24 11140.846016
Rwneg115_25 in115 sn25 3183.098862
Rwneg115_26 in115 sn26 11140.846016
Rwneg115_27 in115 sn27 3183.098862
Rwneg115_28 in115 sn28 11140.846016
Rwneg115_29 in115 sn29 11140.846016
Rwneg115_30 in115 sn30 11140.846016
Rwneg115_31 in115 sn31 11140.846016
Rwneg115_32 in115 sn32 11140.846016
Rwneg115_33 in115 sn33 11140.846016
Rwneg115_34 in115 sn34 11140.846016
Rwneg115_35 in115 sn35 11140.846016
Rwneg115_36 in115 sn36 11140.846016
Rwneg115_37 in115 sn37 11140.846016
Rwneg115_38 in115 sn38 11140.846016
Rwneg115_39 in115 sn39 3183.098862
Rwneg115_40 in115 sn40 11140.846016
Rwneg115_41 in115 sn41 3183.098862
Rwneg115_42 in115 sn42 11140.846016
Rwneg115_43 in115 sn43 3183.098862
Rwneg115_44 in115 sn44 11140.846016
Rwneg115_45 in115 sn45 3183.098862
Rwneg115_46 in115 sn46 11140.846016
Rwneg115_47 in115 sn47 11140.846016
Rwneg115_48 in115 sn48 11140.846016
Rwneg115_49 in115 sn49 11140.846016
Rwneg115_50 in115 sn50 11140.846016
Rwneg115_51 in115 sn51 11140.846016
Rwneg115_52 in115 sn52 3183.098862
Rwneg115_53 in115 sn53 11140.846016
Rwneg115_54 in115 sn54 11140.846016
Rwneg115_55 in115 sn55 3183.098862
Rwneg115_56 in115 sn56 11140.846016
Rwneg115_57 in115 sn57 3183.098862
Rwneg115_58 in115 sn58 11140.846016
Rwneg115_59 in115 sn59 3183.098862
Rwneg115_60 in115 sn60 3183.098862
Rwneg115_61 in115 sn61 3183.098862
Rwneg115_62 in115 sn62 11140.846016
Rwneg115_63 in115 sn63 11140.846016
Rwneg115_64 in115 sn64 11140.846016
Rwneg115_65 in115 sn65 3183.098862
Rwneg115_66 in115 sn66 11140.846016
Rwneg115_67 in115 sn67 11140.846016
Rwneg115_68 in115 sn68 11140.846016
Rwneg115_69 in115 sn69 11140.846016
Rwneg115_70 in115 sn70 11140.846016
Rwneg115_71 in115 sn71 3183.098862
Rwneg115_72 in115 sn72 11140.846016
Rwneg115_73 in115 sn73 11140.846016
Rwneg115_74 in115 sn74 11140.846016
Rwneg115_75 in115 sn75 3183.098862
Rwneg115_76 in115 sn76 11140.846016
Rwneg115_77 in115 sn77 3183.098862
Rwneg115_78 in115 sn78 11140.846016
Rwneg115_79 in115 sn79 3183.098862
Rwneg115_80 in115 sn80 3183.098862
Rwneg115_81 in115 sn81 3183.098862
Rwneg115_82 in115 sn82 11140.846016
Rwneg115_83 in115 sn83 11140.846016
Rwneg115_84 in115 sn84 11140.846016
Rwneg115_85 in115 sn85 11140.846016
Rwneg115_86 in115 sn86 11140.846016
Rwneg115_87 in115 sn87 3183.098862
Rwneg115_88 in115 sn88 11140.846016
Rwneg115_89 in115 sn89 3183.098862
Rwneg115_90 in115 sn90 11140.846016
Rwneg115_91 in115 sn91 3183.098862
Rwneg115_92 in115 sn92 11140.846016
Rwneg115_93 in115 sn93 11140.846016
Rwneg115_94 in115 sn94 11140.846016
Rwneg115_95 in115 sn95 11140.846016
Rwneg115_96 in115 sn96 11140.846016
Rwneg115_97 in115 sn97 11140.846016
Rwneg115_98 in115 sn98 11140.846016
Rwneg115_99 in115 sn99 3183.098862
Rwneg115_100 in115 sn100 11140.846016
Rwneg116_1 in116 sn1 3183.098862
Rwneg116_2 in116 sn2 3183.098862
Rwneg116_3 in116 sn3 11140.846016
Rwneg116_4 in116 sn4 3183.098862
Rwneg116_5 in116 sn5 3183.098862
Rwneg116_6 in116 sn6 11140.846016
Rwneg116_7 in116 sn7 3183.098862
Rwneg116_8 in116 sn8 3183.098862
Rwneg116_9 in116 sn9 11140.846016
Rwneg116_10 in116 sn10 11140.846016
Rwneg116_11 in116 sn11 11140.846016
Rwneg116_12 in116 sn12 11140.846016
Rwneg116_13 in116 sn13 11140.846016
Rwneg116_14 in116 sn14 11140.846016
Rwneg116_15 in116 sn15 11140.846016
Rwneg116_16 in116 sn16 11140.846016
Rwneg116_17 in116 sn17 11140.846016
Rwneg116_18 in116 sn18 11140.846016
Rwneg116_19 in116 sn19 11140.846016
Rwneg116_20 in116 sn20 11140.846016
Rwneg116_21 in116 sn21 11140.846016
Rwneg116_22 in116 sn22 11140.846016
Rwneg116_23 in116 sn23 3183.098862
Rwneg116_24 in116 sn24 11140.846016
Rwneg116_25 in116 sn25 3183.098862
Rwneg116_26 in116 sn26 3183.098862
Rwneg116_27 in116 sn27 11140.846016
Rwneg116_28 in116 sn28 3183.098862
Rwneg116_29 in116 sn29 3183.098862
Rwneg116_30 in116 sn30 11140.846016
Rwneg116_31 in116 sn31 3183.098862
Rwneg116_32 in116 sn32 3183.098862
Rwneg116_33 in116 sn33 11140.846016
Rwneg116_34 in116 sn34 3183.098862
Rwneg116_35 in116 sn35 11140.846016
Rwneg116_36 in116 sn36 3183.098862
Rwneg116_37 in116 sn37 11140.846016
Rwneg116_38 in116 sn38 11140.846016
Rwneg116_39 in116 sn39 3183.098862
Rwneg116_40 in116 sn40 3183.098862
Rwneg116_41 in116 sn41 11140.846016
Rwneg116_42 in116 sn42 11140.846016
Rwneg116_43 in116 sn43 11140.846016
Rwneg116_44 in116 sn44 11140.846016
Rwneg116_45 in116 sn45 11140.846016
Rwneg116_46 in116 sn46 11140.846016
Rwneg116_47 in116 sn47 3183.098862
Rwneg116_48 in116 sn48 11140.846016
Rwneg116_49 in116 sn49 3183.098862
Rwneg116_50 in116 sn50 11140.846016
Rwneg116_51 in116 sn51 3183.098862
Rwneg116_52 in116 sn52 3183.098862
Rwneg116_53 in116 sn53 11140.846016
Rwneg116_54 in116 sn54 11140.846016
Rwneg116_55 in116 sn55 11140.846016
Rwneg116_56 in116 sn56 3183.098862
Rwneg116_57 in116 sn57 11140.846016
Rwneg116_58 in116 sn58 3183.098862
Rwneg116_59 in116 sn59 11140.846016
Rwneg116_60 in116 sn60 3183.098862
Rwneg116_61 in116 sn61 3183.098862
Rwneg116_62 in116 sn62 3183.098862
Rwneg116_63 in116 sn63 11140.846016
Rwneg116_64 in116 sn64 11140.846016
Rwneg116_65 in116 sn65 11140.846016
Rwneg116_66 in116 sn66 11140.846016
Rwneg116_67 in116 sn67 3183.098862
Rwneg116_68 in116 sn68 3183.098862
Rwneg116_69 in116 sn69 3183.098862
Rwneg116_70 in116 sn70 3183.098862
Rwneg116_71 in116 sn71 11140.846016
Rwneg116_72 in116 sn72 11140.846016
Rwneg116_73 in116 sn73 11140.846016
Rwneg116_74 in116 sn74 11140.846016
Rwneg116_75 in116 sn75 11140.846016
Rwneg116_76 in116 sn76 11140.846016
Rwneg116_77 in116 sn77 11140.846016
Rwneg116_78 in116 sn78 3183.098862
Rwneg116_79 in116 sn79 11140.846016
Rwneg116_80 in116 sn80 3183.098862
Rwneg116_81 in116 sn81 11140.846016
Rwneg116_82 in116 sn82 11140.846016
Rwneg116_83 in116 sn83 3183.098862
Rwneg116_84 in116 sn84 3183.098862
Rwneg116_85 in116 sn85 11140.846016
Rwneg116_86 in116 sn86 3183.098862
Rwneg116_87 in116 sn87 11140.846016
Rwneg116_88 in116 sn88 11140.846016
Rwneg116_89 in116 sn89 11140.846016
Rwneg116_90 in116 sn90 11140.846016
Rwneg116_91 in116 sn91 11140.846016
Rwneg116_92 in116 sn92 3183.098862
Rwneg116_93 in116 sn93 11140.846016
Rwneg116_94 in116 sn94 3183.098862
Rwneg116_95 in116 sn95 11140.846016
Rwneg116_96 in116 sn96 11140.846016
Rwneg116_97 in116 sn97 3183.098862
Rwneg116_98 in116 sn98 3183.098862
Rwneg116_99 in116 sn99 11140.846016
Rwneg116_100 in116 sn100 11140.846016
Rwneg117_1 in117 sn1 11140.846016
Rwneg117_2 in117 sn2 3183.098862
Rwneg117_3 in117 sn3 3183.098862
Rwneg117_4 in117 sn4 3183.098862
Rwneg117_5 in117 sn5 3183.098862
Rwneg117_6 in117 sn6 3183.098862
Rwneg117_7 in117 sn7 11140.846016
Rwneg117_8 in117 sn8 11140.846016
Rwneg117_9 in117 sn9 3183.098862
Rwneg117_10 in117 sn10 3183.098862
Rwneg117_11 in117 sn11 11140.846016
Rwneg117_12 in117 sn12 3183.098862
Rwneg117_13 in117 sn13 11140.846016
Rwneg117_14 in117 sn14 3183.098862
Rwneg117_15 in117 sn15 11140.846016
Rwneg117_16 in117 sn16 3183.098862
Rwneg117_17 in117 sn17 11140.846016
Rwneg117_18 in117 sn18 3183.098862
Rwneg117_19 in117 sn19 11140.846016
Rwneg117_20 in117 sn20 3183.098862
Rwneg117_21 in117 sn21 11140.846016
Rwneg117_22 in117 sn22 11140.846016
Rwneg117_23 in117 sn23 11140.846016
Rwneg117_24 in117 sn24 3183.098862
Rwneg117_25 in117 sn25 3183.098862
Rwneg117_26 in117 sn26 3183.098862
Rwneg117_27 in117 sn27 11140.846016
Rwneg117_28 in117 sn28 11140.846016
Rwneg117_29 in117 sn29 11140.846016
Rwneg117_30 in117 sn30 11140.846016
Rwneg117_31 in117 sn31 3183.098862
Rwneg117_32 in117 sn32 3183.098862
Rwneg117_33 in117 sn33 3183.098862
Rwneg117_34 in117 sn34 11140.846016
Rwneg117_35 in117 sn35 11140.846016
Rwneg117_36 in117 sn36 11140.846016
Rwneg117_37 in117 sn37 11140.846016
Rwneg117_38 in117 sn38 11140.846016
Rwneg117_39 in117 sn39 3183.098862
Rwneg117_40 in117 sn40 11140.846016
Rwneg117_41 in117 sn41 11140.846016
Rwneg117_42 in117 sn42 3183.098862
Rwneg117_43 in117 sn43 11140.846016
Rwneg117_44 in117 sn44 3183.098862
Rwneg117_45 in117 sn45 3183.098862
Rwneg117_46 in117 sn46 3183.098862
Rwneg117_47 in117 sn47 11140.846016
Rwneg117_48 in117 sn48 3183.098862
Rwneg117_49 in117 sn49 3183.098862
Rwneg117_50 in117 sn50 11140.846016
Rwneg117_51 in117 sn51 11140.846016
Rwneg117_52 in117 sn52 3183.098862
Rwneg117_53 in117 sn53 11140.846016
Rwneg117_54 in117 sn54 11140.846016
Rwneg117_55 in117 sn55 3183.098862
Rwneg117_56 in117 sn56 11140.846016
Rwneg117_57 in117 sn57 11140.846016
Rwneg117_58 in117 sn58 3183.098862
Rwneg117_59 in117 sn59 3183.098862
Rwneg117_60 in117 sn60 3183.098862
Rwneg117_61 in117 sn61 11140.846016
Rwneg117_62 in117 sn62 11140.846016
Rwneg117_63 in117 sn63 11140.846016
Rwneg117_64 in117 sn64 3183.098862
Rwneg117_65 in117 sn65 3183.098862
Rwneg117_66 in117 sn66 3183.098862
Rwneg117_67 in117 sn67 11140.846016
Rwneg117_68 in117 sn68 3183.098862
Rwneg117_69 in117 sn69 3183.098862
Rwneg117_70 in117 sn70 11140.846016
Rwneg117_71 in117 sn71 11140.846016
Rwneg117_72 in117 sn72 3183.098862
Rwneg117_73 in117 sn73 11140.846016
Rwneg117_74 in117 sn74 3183.098862
Rwneg117_75 in117 sn75 11140.846016
Rwneg117_76 in117 sn76 3183.098862
Rwneg117_77 in117 sn77 3183.098862
Rwneg117_78 in117 sn78 3183.098862
Rwneg117_79 in117 sn79 11140.846016
Rwneg117_80 in117 sn80 3183.098862
Rwneg117_81 in117 sn81 11140.846016
Rwneg117_82 in117 sn82 11140.846016
Rwneg117_83 in117 sn83 3183.098862
Rwneg117_84 in117 sn84 3183.098862
Rwneg117_85 in117 sn85 11140.846016
Rwneg117_86 in117 sn86 11140.846016
Rwneg117_87 in117 sn87 11140.846016
Rwneg117_88 in117 sn88 11140.846016
Rwneg117_89 in117 sn89 3183.098862
Rwneg117_90 in117 sn90 11140.846016
Rwneg117_91 in117 sn91 3183.098862
Rwneg117_92 in117 sn92 3183.098862
Rwneg117_93 in117 sn93 3183.098862
Rwneg117_94 in117 sn94 11140.846016
Rwneg117_95 in117 sn95 3183.098862
Rwneg117_96 in117 sn96 3183.098862
Rwneg117_97 in117 sn97 11140.846016
Rwneg117_98 in117 sn98 11140.846016
Rwneg117_99 in117 sn99 3183.098862
Rwneg117_100 in117 sn100 3183.098862
Rwneg118_1 in118 sn1 11140.846016
Rwneg118_2 in118 sn2 11140.846016
Rwneg118_3 in118 sn3 3183.098862
Rwneg118_4 in118 sn4 11140.846016
Rwneg118_5 in118 sn5 3183.098862
Rwneg118_6 in118 sn6 11140.846016
Rwneg118_7 in118 sn7 3183.098862
Rwneg118_8 in118 sn8 3183.098862
Rwneg118_9 in118 sn9 3183.098862
Rwneg118_10 in118 sn10 11140.846016
Rwneg118_11 in118 sn11 11140.846016
Rwneg118_12 in118 sn12 3183.098862
Rwneg118_13 in118 sn13 3183.098862
Rwneg118_14 in118 sn14 11140.846016
Rwneg118_15 in118 sn15 11140.846016
Rwneg118_16 in118 sn16 11140.846016
Rwneg118_17 in118 sn17 3183.098862
Rwneg118_18 in118 sn18 11140.846016
Rwneg118_19 in118 sn19 11140.846016
Rwneg118_20 in118 sn20 11140.846016
Rwneg118_21 in118 sn21 11140.846016
Rwneg118_22 in118 sn22 3183.098862
Rwneg118_23 in118 sn23 3183.098862
Rwneg118_24 in118 sn24 3183.098862
Rwneg118_25 in118 sn25 3183.098862
Rwneg118_26 in118 sn26 3183.098862
Rwneg118_27 in118 sn27 11140.846016
Rwneg118_28 in118 sn28 11140.846016
Rwneg118_29 in118 sn29 11140.846016
Rwneg118_30 in118 sn30 11140.846016
Rwneg118_31 in118 sn31 11140.846016
Rwneg118_32 in118 sn32 3183.098862
Rwneg118_33 in118 sn33 11140.846016
Rwneg118_34 in118 sn34 3183.098862
Rwneg118_35 in118 sn35 3183.098862
Rwneg118_36 in118 sn36 11140.846016
Rwneg118_37 in118 sn37 11140.846016
Rwneg118_38 in118 sn38 11140.846016
Rwneg118_39 in118 sn39 3183.098862
Rwneg118_40 in118 sn40 11140.846016
Rwneg118_41 in118 sn41 11140.846016
Rwneg118_42 in118 sn42 3183.098862
Rwneg118_43 in118 sn43 3183.098862
Rwneg118_44 in118 sn44 11140.846016
Rwneg118_45 in118 sn45 11140.846016
Rwneg118_46 in118 sn46 11140.846016
Rwneg118_47 in118 sn47 11140.846016
Rwneg118_48 in118 sn48 3183.098862
Rwneg118_49 in118 sn49 3183.098862
Rwneg118_50 in118 sn50 11140.846016
Rwneg118_51 in118 sn51 3183.098862
Rwneg118_52 in118 sn52 11140.846016
Rwneg118_53 in118 sn53 11140.846016
Rwneg118_54 in118 sn54 3183.098862
Rwneg118_55 in118 sn55 3183.098862
Rwneg118_56 in118 sn56 11140.846016
Rwneg118_57 in118 sn57 3183.098862
Rwneg118_58 in118 sn58 11140.846016
Rwneg118_59 in118 sn59 3183.098862
Rwneg118_60 in118 sn60 3183.098862
Rwneg118_61 in118 sn61 3183.098862
Rwneg118_62 in118 sn62 3183.098862
Rwneg118_63 in118 sn63 3183.098862
Rwneg118_64 in118 sn64 3183.098862
Rwneg118_65 in118 sn65 11140.846016
Rwneg118_66 in118 sn66 3183.098862
Rwneg118_67 in118 sn67 11140.846016
Rwneg118_68 in118 sn68 3183.098862
Rwneg118_69 in118 sn69 3183.098862
Rwneg118_70 in118 sn70 3183.098862
Rwneg118_71 in118 sn71 11140.846016
Rwneg118_72 in118 sn72 11140.846016
Rwneg118_73 in118 sn73 11140.846016
Rwneg118_74 in118 sn74 11140.846016
Rwneg118_75 in118 sn75 11140.846016
Rwneg118_76 in118 sn76 3183.098862
Rwneg118_77 in118 sn77 3183.098862
Rwneg118_78 in118 sn78 3183.098862
Rwneg118_79 in118 sn79 11140.846016
Rwneg118_80 in118 sn80 3183.098862
Rwneg118_81 in118 sn81 11140.846016
Rwneg118_82 in118 sn82 11140.846016
Rwneg118_83 in118 sn83 11140.846016
Rwneg118_84 in118 sn84 3183.098862
Rwneg118_85 in118 sn85 3183.098862
Rwneg118_86 in118 sn86 3183.098862
Rwneg118_87 in118 sn87 3183.098862
Rwneg118_88 in118 sn88 11140.846016
Rwneg118_89 in118 sn89 3183.098862
Rwneg118_90 in118 sn90 11140.846016
Rwneg118_91 in118 sn91 11140.846016
Rwneg118_92 in118 sn92 3183.098862
Rwneg118_93 in118 sn93 11140.846016
Rwneg118_94 in118 sn94 11140.846016
Rwneg118_95 in118 sn95 3183.098862
Rwneg118_96 in118 sn96 11140.846016
Rwneg118_97 in118 sn97 3183.098862
Rwneg118_98 in118 sn98 3183.098862
Rwneg118_99 in118 sn99 3183.098862
Rwneg118_100 in118 sn100 3183.098862
Rwneg119_1 in119 sn1 11140.846016
Rwneg119_2 in119 sn2 11140.846016
Rwneg119_3 in119 sn3 3183.098862
Rwneg119_4 in119 sn4 3183.098862
Rwneg119_5 in119 sn5 11140.846016
Rwneg119_6 in119 sn6 3183.098862
Rwneg119_7 in119 sn7 3183.098862
Rwneg119_8 in119 sn8 11140.846016
Rwneg119_9 in119 sn9 3183.098862
Rwneg119_10 in119 sn10 11140.846016
Rwneg119_11 in119 sn11 3183.098862
Rwneg119_12 in119 sn12 11140.846016
Rwneg119_13 in119 sn13 3183.098862
Rwneg119_14 in119 sn14 11140.846016
Rwneg119_15 in119 sn15 11140.846016
Rwneg119_16 in119 sn16 11140.846016
Rwneg119_17 in119 sn17 11140.846016
Rwneg119_18 in119 sn18 3183.098862
Rwneg119_19 in119 sn19 3183.098862
Rwneg119_20 in119 sn20 11140.846016
Rwneg119_21 in119 sn21 11140.846016
Rwneg119_22 in119 sn22 3183.098862
Rwneg119_23 in119 sn23 3183.098862
Rwneg119_24 in119 sn24 11140.846016
Rwneg119_25 in119 sn25 3183.098862
Rwneg119_26 in119 sn26 11140.846016
Rwneg119_27 in119 sn27 11140.846016
Rwneg119_28 in119 sn28 3183.098862
Rwneg119_29 in119 sn29 11140.846016
Rwneg119_30 in119 sn30 11140.846016
Rwneg119_31 in119 sn31 3183.098862
Rwneg119_32 in119 sn32 11140.846016
Rwneg119_33 in119 sn33 11140.846016
Rwneg119_34 in119 sn34 11140.846016
Rwneg119_35 in119 sn35 11140.846016
Rwneg119_36 in119 sn36 11140.846016
Rwneg119_37 in119 sn37 3183.098862
Rwneg119_38 in119 sn38 11140.846016
Rwneg119_39 in119 sn39 11140.846016
Rwneg119_40 in119 sn40 11140.846016
Rwneg119_41 in119 sn41 3183.098862
Rwneg119_42 in119 sn42 11140.846016
Rwneg119_43 in119 sn43 3183.098862
Rwneg119_44 in119 sn44 11140.846016
Rwneg119_45 in119 sn45 3183.098862
Rwneg119_46 in119 sn46 11140.846016
Rwneg119_47 in119 sn47 11140.846016
Rwneg119_48 in119 sn48 11140.846016
Rwneg119_49 in119 sn49 11140.846016
Rwneg119_50 in119 sn50 11140.846016
Rwneg119_51 in119 sn51 11140.846016
Rwneg119_52 in119 sn52 11140.846016
Rwneg119_53 in119 sn53 3183.098862
Rwneg119_54 in119 sn54 11140.846016
Rwneg119_55 in119 sn55 11140.846016
Rwneg119_56 in119 sn56 11140.846016
Rwneg119_57 in119 sn57 3183.098862
Rwneg119_58 in119 sn58 11140.846016
Rwneg119_59 in119 sn59 3183.098862
Rwneg119_60 in119 sn60 3183.098862
Rwneg119_61 in119 sn61 3183.098862
Rwneg119_62 in119 sn62 11140.846016
Rwneg119_63 in119 sn63 11140.846016
Rwneg119_64 in119 sn64 3183.098862
Rwneg119_65 in119 sn65 3183.098862
Rwneg119_66 in119 sn66 11140.846016
Rwneg119_67 in119 sn67 11140.846016
Rwneg119_68 in119 sn68 11140.846016
Rwneg119_69 in119 sn69 11140.846016
Rwneg119_70 in119 sn70 11140.846016
Rwneg119_71 in119 sn71 3183.098862
Rwneg119_72 in119 sn72 3183.098862
Rwneg119_73 in119 sn73 3183.098862
Rwneg119_74 in119 sn74 11140.846016
Rwneg119_75 in119 sn75 3183.098862
Rwneg119_76 in119 sn76 3183.098862
Rwneg119_77 in119 sn77 3183.098862
Rwneg119_78 in119 sn78 3183.098862
Rwneg119_79 in119 sn79 11140.846016
Rwneg119_80 in119 sn80 3183.098862
Rwneg119_81 in119 sn81 3183.098862
Rwneg119_82 in119 sn82 11140.846016
Rwneg119_83 in119 sn83 3183.098862
Rwneg119_84 in119 sn84 3183.098862
Rwneg119_85 in119 sn85 11140.846016
Rwneg119_86 in119 sn86 3183.098862
Rwneg119_87 in119 sn87 11140.846016
Rwneg119_88 in119 sn88 11140.846016
Rwneg119_89 in119 sn89 3183.098862
Rwneg119_90 in119 sn90 11140.846016
Rwneg119_91 in119 sn91 3183.098862
Rwneg119_92 in119 sn92 3183.098862
Rwneg119_93 in119 sn93 3183.098862
Rwneg119_94 in119 sn94 11140.846016
Rwneg119_95 in119 sn95 11140.846016
Rwneg119_96 in119 sn96 3183.098862
Rwneg119_97 in119 sn97 3183.098862
Rwneg119_98 in119 sn98 11140.846016
Rwneg119_99 in119 sn99 11140.846016
Rwneg119_100 in119 sn100 11140.846016
Rwneg120_1 in120 sn1 11140.846016
Rwneg120_2 in120 sn2 11140.846016
Rwneg120_3 in120 sn3 3183.098862
Rwneg120_4 in120 sn4 11140.846016
Rwneg120_5 in120 sn5 3183.098862
Rwneg120_6 in120 sn6 11140.846016
Rwneg120_7 in120 sn7 3183.098862
Rwneg120_8 in120 sn8 11140.846016
Rwneg120_9 in120 sn9 11140.846016
Rwneg120_10 in120 sn10 11140.846016
Rwneg120_11 in120 sn11 11140.846016
Rwneg120_12 in120 sn12 3183.098862
Rwneg120_13 in120 sn13 3183.098862
Rwneg120_14 in120 sn14 11140.846016
Rwneg120_15 in120 sn15 11140.846016
Rwneg120_16 in120 sn16 11140.846016
Rwneg120_17 in120 sn17 11140.846016
Rwneg120_18 in120 sn18 11140.846016
Rwneg120_19 in120 sn19 3183.098862
Rwneg120_20 in120 sn20 11140.846016
Rwneg120_21 in120 sn21 3183.098862
Rwneg120_22 in120 sn22 11140.846016
Rwneg120_23 in120 sn23 3183.098862
Rwneg120_24 in120 sn24 3183.098862
Rwneg120_25 in120 sn25 3183.098862
Rwneg120_26 in120 sn26 11140.846016
Rwneg120_27 in120 sn27 11140.846016
Rwneg120_28 in120 sn28 3183.098862
Rwneg120_29 in120 sn29 11140.846016
Rwneg120_30 in120 sn30 11140.846016
Rwneg120_31 in120 sn31 11140.846016
Rwneg120_32 in120 sn32 11140.846016
Rwneg120_33 in120 sn33 11140.846016
Rwneg120_34 in120 sn34 11140.846016
Rwneg120_35 in120 sn35 3183.098862
Rwneg120_36 in120 sn36 11140.846016
Rwneg120_37 in120 sn37 3183.098862
Rwneg120_38 in120 sn38 11140.846016
Rwneg120_39 in120 sn39 3183.098862
Rwneg120_40 in120 sn40 3183.098862
Rwneg120_41 in120 sn41 3183.098862
Rwneg120_42 in120 sn42 3183.098862
Rwneg120_43 in120 sn43 11140.846016
Rwneg120_44 in120 sn44 11140.846016
Rwneg120_45 in120 sn45 11140.846016
Rwneg120_46 in120 sn46 11140.846016
Rwneg120_47 in120 sn47 11140.846016
Rwneg120_48 in120 sn48 11140.846016
Rwneg120_49 in120 sn49 11140.846016
Rwneg120_50 in120 sn50 11140.846016
Rwneg120_51 in120 sn51 3183.098862
Rwneg120_52 in120 sn52 3183.098862
Rwneg120_53 in120 sn53 11140.846016
Rwneg120_54 in120 sn54 11140.846016
Rwneg120_55 in120 sn55 11140.846016
Rwneg120_56 in120 sn56 11140.846016
Rwneg120_57 in120 sn57 3183.098862
Rwneg120_58 in120 sn58 11140.846016
Rwneg120_59 in120 sn59 3183.098862
Rwneg120_60 in120 sn60 11140.846016
Rwneg120_61 in120 sn61 11140.846016
Rwneg120_62 in120 sn62 3183.098862
Rwneg120_63 in120 sn63 11140.846016
Rwneg120_64 in120 sn64 11140.846016
Rwneg120_65 in120 sn65 11140.846016
Rwneg120_66 in120 sn66 3183.098862
Rwneg120_67 in120 sn67 11140.846016
Rwneg120_68 in120 sn68 11140.846016
Rwneg120_69 in120 sn69 11140.846016
Rwneg120_70 in120 sn70 11140.846016
Rwneg120_71 in120 sn71 3183.098862
Rwneg120_72 in120 sn72 3183.098862
Rwneg120_73 in120 sn73 3183.098862
Rwneg120_74 in120 sn74 3183.098862
Rwneg120_75 in120 sn75 3183.098862
Rwneg120_76 in120 sn76 11140.846016
Rwneg120_77 in120 sn77 3183.098862
Rwneg120_78 in120 sn78 11140.846016
Rwneg120_79 in120 sn79 3183.098862
Rwneg120_80 in120 sn80 3183.098862
Rwneg120_81 in120 sn81 3183.098862
Rwneg120_82 in120 sn82 11140.846016
Rwneg120_83 in120 sn83 3183.098862
Rwneg120_84 in120 sn84 3183.098862
Rwneg120_85 in120 sn85 11140.846016
Rwneg120_86 in120 sn86 3183.098862
Rwneg120_87 in120 sn87 11140.846016
Rwneg120_88 in120 sn88 3183.098862
Rwneg120_89 in120 sn89 3183.098862
Rwneg120_90 in120 sn90 11140.846016
Rwneg120_91 in120 sn91 11140.846016
Rwneg120_92 in120 sn92 3183.098862
Rwneg120_93 in120 sn93 11140.846016
Rwneg120_94 in120 sn94 11140.846016
Rwneg120_95 in120 sn95 3183.098862
Rwneg120_96 in120 sn96 11140.846016
Rwneg120_97 in120 sn97 11140.846016
Rwneg120_98 in120 sn98 3183.098862
Rwneg120_99 in120 sn99 3183.098862
Rwneg120_100 in120 sn100 11140.846016
Rwneg121_1 in121 sn1 3183.098862
Rwneg121_2 in121 sn2 3183.098862
Rwneg121_3 in121 sn3 11140.846016
Rwneg121_4 in121 sn4 11140.846016
Rwneg121_5 in121 sn5 3183.098862
Rwneg121_6 in121 sn6 11140.846016
Rwneg121_7 in121 sn7 3183.098862
Rwneg121_8 in121 sn8 11140.846016
Rwneg121_9 in121 sn9 11140.846016
Rwneg121_10 in121 sn10 11140.846016
Rwneg121_11 in121 sn11 11140.846016
Rwneg121_12 in121 sn12 3183.098862
Rwneg121_13 in121 sn13 11140.846016
Rwneg121_14 in121 sn14 3183.098862
Rwneg121_15 in121 sn15 11140.846016
Rwneg121_16 in121 sn16 3183.098862
Rwneg121_17 in121 sn17 3183.098862
Rwneg121_18 in121 sn18 3183.098862
Rwneg121_19 in121 sn19 11140.846016
Rwneg121_20 in121 sn20 11140.846016
Rwneg121_21 in121 sn21 11140.846016
Rwneg121_22 in121 sn22 11140.846016
Rwneg121_23 in121 sn23 3183.098862
Rwneg121_24 in121 sn24 11140.846016
Rwneg121_25 in121 sn25 3183.098862
Rwneg121_26 in121 sn26 3183.098862
Rwneg121_27 in121 sn27 3183.098862
Rwneg121_28 in121 sn28 3183.098862
Rwneg121_29 in121 sn29 3183.098862
Rwneg121_30 in121 sn30 3183.098862
Rwneg121_31 in121 sn31 11140.846016
Rwneg121_32 in121 sn32 3183.098862
Rwneg121_33 in121 sn33 11140.846016
Rwneg121_34 in121 sn34 3183.098862
Rwneg121_35 in121 sn35 11140.846016
Rwneg121_36 in121 sn36 11140.846016
Rwneg121_37 in121 sn37 11140.846016
Rwneg121_38 in121 sn38 3183.098862
Rwneg121_39 in121 sn39 11140.846016
Rwneg121_40 in121 sn40 11140.846016
Rwneg121_41 in121 sn41 11140.846016
Rwneg121_42 in121 sn42 3183.098862
Rwneg121_43 in121 sn43 11140.846016
Rwneg121_44 in121 sn44 3183.098862
Rwneg121_45 in121 sn45 3183.098862
Rwneg121_46 in121 sn46 3183.098862
Rwneg121_47 in121 sn47 3183.098862
Rwneg121_48 in121 sn48 3183.098862
Rwneg121_49 in121 sn49 11140.846016
Rwneg121_50 in121 sn50 3183.098862
Rwneg121_51 in121 sn51 3183.098862
Rwneg121_52 in121 sn52 11140.846016
Rwneg121_53 in121 sn53 3183.098862
Rwneg121_54 in121 sn54 11140.846016
Rwneg121_55 in121 sn55 3183.098862
Rwneg121_56 in121 sn56 11140.846016
Rwneg121_57 in121 sn57 3183.098862
Rwneg121_58 in121 sn58 11140.846016
Rwneg121_59 in121 sn59 3183.098862
Rwneg121_60 in121 sn60 11140.846016
Rwneg121_61 in121 sn61 3183.098862
Rwneg121_62 in121 sn62 3183.098862
Rwneg121_63 in121 sn63 3183.098862
Rwneg121_64 in121 sn64 3183.098862
Rwneg121_65 in121 sn65 11140.846016
Rwneg121_66 in121 sn66 3183.098862
Rwneg121_67 in121 sn67 11140.846016
Rwneg121_68 in121 sn68 11140.846016
Rwneg121_69 in121 sn69 3183.098862
Rwneg121_70 in121 sn70 11140.846016
Rwneg121_71 in121 sn71 11140.846016
Rwneg121_72 in121 sn72 11140.846016
Rwneg121_73 in121 sn73 11140.846016
Rwneg121_74 in121 sn74 11140.846016
Rwneg121_75 in121 sn75 11140.846016
Rwneg121_76 in121 sn76 3183.098862
Rwneg121_77 in121 sn77 3183.098862
Rwneg121_78 in121 sn78 11140.846016
Rwneg121_79 in121 sn79 11140.846016
Rwneg121_80 in121 sn80 3183.098862
Rwneg121_81 in121 sn81 3183.098862
Rwneg121_82 in121 sn82 3183.098862
Rwneg121_83 in121 sn83 11140.846016
Rwneg121_84 in121 sn84 11140.846016
Rwneg121_85 in121 sn85 11140.846016
Rwneg121_86 in121 sn86 3183.098862
Rwneg121_87 in121 sn87 3183.098862
Rwneg121_88 in121 sn88 3183.098862
Rwneg121_89 in121 sn89 11140.846016
Rwneg121_90 in121 sn90 11140.846016
Rwneg121_91 in121 sn91 11140.846016
Rwneg121_92 in121 sn92 11140.846016
Rwneg121_93 in121 sn93 11140.846016
Rwneg121_94 in121 sn94 3183.098862
Rwneg121_95 in121 sn95 11140.846016
Rwneg121_96 in121 sn96 11140.846016
Rwneg121_97 in121 sn97 11140.846016
Rwneg121_98 in121 sn98 11140.846016
Rwneg121_99 in121 sn99 11140.846016
Rwneg121_100 in121 sn100 3183.098862
Rwneg122_1 in122 sn1 11140.846016
Rwneg122_2 in122 sn2 3183.098862
Rwneg122_3 in122 sn3 3183.098862
Rwneg122_4 in122 sn4 11140.846016
Rwneg122_5 in122 sn5 11140.846016
Rwneg122_6 in122 sn6 3183.098862
Rwneg122_7 in122 sn7 3183.098862
Rwneg122_8 in122 sn8 11140.846016
Rwneg122_9 in122 sn9 11140.846016
Rwneg122_10 in122 sn10 3183.098862
Rwneg122_11 in122 sn11 3183.098862
Rwneg122_12 in122 sn12 3183.098862
Rwneg122_13 in122 sn13 11140.846016
Rwneg122_14 in122 sn14 3183.098862
Rwneg122_15 in122 sn15 11140.846016
Rwneg122_16 in122 sn16 3183.098862
Rwneg122_17 in122 sn17 11140.846016
Rwneg122_18 in122 sn18 3183.098862
Rwneg122_19 in122 sn19 11140.846016
Rwneg122_20 in122 sn20 11140.846016
Rwneg122_21 in122 sn21 3183.098862
Rwneg122_22 in122 sn22 11140.846016
Rwneg122_23 in122 sn23 3183.098862
Rwneg122_24 in122 sn24 3183.098862
Rwneg122_25 in122 sn25 3183.098862
Rwneg122_26 in122 sn26 3183.098862
Rwneg122_27 in122 sn27 11140.846016
Rwneg122_28 in122 sn28 11140.846016
Rwneg122_29 in122 sn29 3183.098862
Rwneg122_30 in122 sn30 3183.098862
Rwneg122_31 in122 sn31 3183.098862
Rwneg122_32 in122 sn32 11140.846016
Rwneg122_33 in122 sn33 11140.846016
Rwneg122_34 in122 sn34 3183.098862
Rwneg122_35 in122 sn35 11140.846016
Rwneg122_36 in122 sn36 11140.846016
Rwneg122_37 in122 sn37 11140.846016
Rwneg122_38 in122 sn38 3183.098862
Rwneg122_39 in122 sn39 3183.098862
Rwneg122_40 in122 sn40 11140.846016
Rwneg122_41 in122 sn41 11140.846016
Rwneg122_42 in122 sn42 3183.098862
Rwneg122_43 in122 sn43 11140.846016
Rwneg122_44 in122 sn44 11140.846016
Rwneg122_45 in122 sn45 3183.098862
Rwneg122_46 in122 sn46 3183.098862
Rwneg122_47 in122 sn47 3183.098862
Rwneg122_48 in122 sn48 11140.846016
Rwneg122_49 in122 sn49 11140.846016
Rwneg122_50 in122 sn50 11140.846016
Rwneg122_51 in122 sn51 3183.098862
Rwneg122_52 in122 sn52 11140.846016
Rwneg122_53 in122 sn53 3183.098862
Rwneg122_54 in122 sn54 3183.098862
Rwneg122_55 in122 sn55 11140.846016
Rwneg122_56 in122 sn56 11140.846016
Rwneg122_57 in122 sn57 3183.098862
Rwneg122_58 in122 sn58 3183.098862
Rwneg122_59 in122 sn59 11140.846016
Rwneg122_60 in122 sn60 3183.098862
Rwneg122_61 in122 sn61 11140.846016
Rwneg122_62 in122 sn62 3183.098862
Rwneg122_63 in122 sn63 11140.846016
Rwneg122_64 in122 sn64 3183.098862
Rwneg122_65 in122 sn65 3183.098862
Rwneg122_66 in122 sn66 11140.846016
Rwneg122_67 in122 sn67 11140.846016
Rwneg122_68 in122 sn68 3183.098862
Rwneg122_69 in122 sn69 3183.098862
Rwneg122_70 in122 sn70 11140.846016
Rwneg122_71 in122 sn71 3183.098862
Rwneg122_72 in122 sn72 11140.846016
Rwneg122_73 in122 sn73 11140.846016
Rwneg122_74 in122 sn74 3183.098862
Rwneg122_75 in122 sn75 11140.846016
Rwneg122_76 in122 sn76 11140.846016
Rwneg122_77 in122 sn77 3183.098862
Rwneg122_78 in122 sn78 11140.846016
Rwneg122_79 in122 sn79 11140.846016
Rwneg122_80 in122 sn80 3183.098862
Rwneg122_81 in122 sn81 11140.846016
Rwneg122_82 in122 sn82 11140.846016
Rwneg122_83 in122 sn83 3183.098862
Rwneg122_84 in122 sn84 11140.846016
Rwneg122_85 in122 sn85 11140.846016
Rwneg122_86 in122 sn86 3183.098862
Rwneg122_87 in122 sn87 11140.846016
Rwneg122_88 in122 sn88 3183.098862
Rwneg122_89 in122 sn89 3183.098862
Rwneg122_90 in122 sn90 3183.098862
Rwneg122_91 in122 sn91 11140.846016
Rwneg122_92 in122 sn92 11140.846016
Rwneg122_93 in122 sn93 11140.846016
Rwneg122_94 in122 sn94 11140.846016
Rwneg122_95 in122 sn95 3183.098862
Rwneg122_96 in122 sn96 3183.098862
Rwneg122_97 in122 sn97 11140.846016
Rwneg122_98 in122 sn98 3183.098862
Rwneg122_99 in122 sn99 3183.098862
Rwneg122_100 in122 sn100 3183.098862
Rwneg123_1 in123 sn1 3183.098862
Rwneg123_2 in123 sn2 3183.098862
Rwneg123_3 in123 sn3 3183.098862
Rwneg123_4 in123 sn4 3183.098862
Rwneg123_5 in123 sn5 3183.098862
Rwneg123_6 in123 sn6 11140.846016
Rwneg123_7 in123 sn7 11140.846016
Rwneg123_8 in123 sn8 3183.098862
Rwneg123_9 in123 sn9 3183.098862
Rwneg123_10 in123 sn10 11140.846016
Rwneg123_11 in123 sn11 3183.098862
Rwneg123_12 in123 sn12 3183.098862
Rwneg123_13 in123 sn13 3183.098862
Rwneg123_14 in123 sn14 11140.846016
Rwneg123_15 in123 sn15 11140.846016
Rwneg123_16 in123 sn16 3183.098862
Rwneg123_17 in123 sn17 3183.098862
Rwneg123_18 in123 sn18 3183.098862
Rwneg123_19 in123 sn19 3183.098862
Rwneg123_20 in123 sn20 3183.098862
Rwneg123_21 in123 sn21 3183.098862
Rwneg123_22 in123 sn22 3183.098862
Rwneg123_23 in123 sn23 3183.098862
Rwneg123_24 in123 sn24 3183.098862
Rwneg123_25 in123 sn25 3183.098862
Rwneg123_26 in123 sn26 11140.846016
Rwneg123_27 in123 sn27 11140.846016
Rwneg123_28 in123 sn28 11140.846016
Rwneg123_29 in123 sn29 11140.846016
Rwneg123_30 in123 sn30 11140.846016
Rwneg123_31 in123 sn31 3183.098862
Rwneg123_32 in123 sn32 11140.846016
Rwneg123_33 in123 sn33 11140.846016
Rwneg123_34 in123 sn34 11140.846016
Rwneg123_35 in123 sn35 11140.846016
Rwneg123_36 in123 sn36 11140.846016
Rwneg123_37 in123 sn37 11140.846016
Rwneg123_38 in123 sn38 3183.098862
Rwneg123_39 in123 sn39 11140.846016
Rwneg123_40 in123 sn40 3183.098862
Rwneg123_41 in123 sn41 11140.846016
Rwneg123_42 in123 sn42 11140.846016
Rwneg123_43 in123 sn43 11140.846016
Rwneg123_44 in123 sn44 11140.846016
Rwneg123_45 in123 sn45 3183.098862
Rwneg123_46 in123 sn46 11140.846016
Rwneg123_47 in123 sn47 3183.098862
Rwneg123_48 in123 sn48 11140.846016
Rwneg123_49 in123 sn49 3183.098862
Rwneg123_50 in123 sn50 3183.098862
Rwneg123_51 in123 sn51 3183.098862
Rwneg123_52 in123 sn52 3183.098862
Rwneg123_53 in123 sn53 11140.846016
Rwneg123_54 in123 sn54 3183.098862
Rwneg123_55 in123 sn55 3183.098862
Rwneg123_56 in123 sn56 11140.846016
Rwneg123_57 in123 sn57 11140.846016
Rwneg123_58 in123 sn58 3183.098862
Rwneg123_59 in123 sn59 3183.098862
Rwneg123_60 in123 sn60 3183.098862
Rwneg123_61 in123 sn61 11140.846016
Rwneg123_62 in123 sn62 11140.846016
Rwneg123_63 in123 sn63 3183.098862
Rwneg123_64 in123 sn64 11140.846016
Rwneg123_65 in123 sn65 3183.098862
Rwneg123_66 in123 sn66 3183.098862
Rwneg123_67 in123 sn67 11140.846016
Rwneg123_68 in123 sn68 3183.098862
Rwneg123_69 in123 sn69 3183.098862
Rwneg123_70 in123 sn70 11140.846016
Rwneg123_71 in123 sn71 11140.846016
Rwneg123_72 in123 sn72 3183.098862
Rwneg123_73 in123 sn73 3183.098862
Rwneg123_74 in123 sn74 3183.098862
Rwneg123_75 in123 sn75 11140.846016
Rwneg123_76 in123 sn76 11140.846016
Rwneg123_77 in123 sn77 11140.846016
Rwneg123_78 in123 sn78 3183.098862
Rwneg123_79 in123 sn79 11140.846016
Rwneg123_80 in123 sn80 11140.846016
Rwneg123_81 in123 sn81 3183.098862
Rwneg123_82 in123 sn82 3183.098862
Rwneg123_83 in123 sn83 3183.098862
Rwneg123_84 in123 sn84 3183.098862
Rwneg123_85 in123 sn85 11140.846016
Rwneg123_86 in123 sn86 3183.098862
Rwneg123_87 in123 sn87 11140.846016
Rwneg123_88 in123 sn88 11140.846016
Rwneg123_89 in123 sn89 11140.846016
Rwneg123_90 in123 sn90 3183.098862
Rwneg123_91 in123 sn91 11140.846016
Rwneg123_92 in123 sn92 3183.098862
Rwneg123_93 in123 sn93 3183.098862
Rwneg123_94 in123 sn94 3183.098862
Rwneg123_95 in123 sn95 11140.846016
Rwneg123_96 in123 sn96 3183.098862
Rwneg123_97 in123 sn97 3183.098862
Rwneg123_98 in123 sn98 3183.098862
Rwneg123_99 in123 sn99 11140.846016
Rwneg123_100 in123 sn100 11140.846016
Rwneg124_1 in124 sn1 3183.098862
Rwneg124_2 in124 sn2 3183.098862
Rwneg124_3 in124 sn3 3183.098862
Rwneg124_4 in124 sn4 3183.098862
Rwneg124_5 in124 sn5 11140.846016
Rwneg124_6 in124 sn6 11140.846016
Rwneg124_7 in124 sn7 3183.098862
Rwneg124_8 in124 sn8 11140.846016
Rwneg124_9 in124 sn9 3183.098862
Rwneg124_10 in124 sn10 3183.098862
Rwneg124_11 in124 sn11 3183.098862
Rwneg124_12 in124 sn12 3183.098862
Rwneg124_13 in124 sn13 3183.098862
Rwneg124_14 in124 sn14 11140.846016
Rwneg124_15 in124 sn15 3183.098862
Rwneg124_16 in124 sn16 11140.846016
Rwneg124_17 in124 sn17 11140.846016
Rwneg124_18 in124 sn18 3183.098862
Rwneg124_19 in124 sn19 11140.846016
Rwneg124_20 in124 sn20 3183.098862
Rwneg124_21 in124 sn21 11140.846016
Rwneg124_22 in124 sn22 11140.846016
Rwneg124_23 in124 sn23 3183.098862
Rwneg124_24 in124 sn24 11140.846016
Rwneg124_25 in124 sn25 11140.846016
Rwneg124_26 in124 sn26 11140.846016
Rwneg124_27 in124 sn27 3183.098862
Rwneg124_28 in124 sn28 11140.846016
Rwneg124_29 in124 sn29 11140.846016
Rwneg124_30 in124 sn30 11140.846016
Rwneg124_31 in124 sn31 11140.846016
Rwneg124_32 in124 sn32 3183.098862
Rwneg124_33 in124 sn33 3183.098862
Rwneg124_34 in124 sn34 11140.846016
Rwneg124_35 in124 sn35 3183.098862
Rwneg124_36 in124 sn36 11140.846016
Rwneg124_37 in124 sn37 3183.098862
Rwneg124_38 in124 sn38 11140.846016
Rwneg124_39 in124 sn39 3183.098862
Rwneg124_40 in124 sn40 3183.098862
Rwneg124_41 in124 sn41 3183.098862
Rwneg124_42 in124 sn42 3183.098862
Rwneg124_43 in124 sn43 3183.098862
Rwneg124_44 in124 sn44 3183.098862
Rwneg124_45 in124 sn45 3183.098862
Rwneg124_46 in124 sn46 3183.098862
Rwneg124_47 in124 sn47 3183.098862
Rwneg124_48 in124 sn48 3183.098862
Rwneg124_49 in124 sn49 3183.098862
Rwneg124_50 in124 sn50 11140.846016
Rwneg124_51 in124 sn51 3183.098862
Rwneg124_52 in124 sn52 3183.098862
Rwneg124_53 in124 sn53 11140.846016
Rwneg124_54 in124 sn54 11140.846016
Rwneg124_55 in124 sn55 11140.846016
Rwneg124_56 in124 sn56 3183.098862
Rwneg124_57 in124 sn57 11140.846016
Rwneg124_58 in124 sn58 11140.846016
Rwneg124_59 in124 sn59 3183.098862
Rwneg124_60 in124 sn60 11140.846016
Rwneg124_61 in124 sn61 3183.098862
Rwneg124_62 in124 sn62 3183.098862
Rwneg124_63 in124 sn63 3183.098862
Rwneg124_64 in124 sn64 3183.098862
Rwneg124_65 in124 sn65 3183.098862
Rwneg124_66 in124 sn66 11140.846016
Rwneg124_67 in124 sn67 11140.846016
Rwneg124_68 in124 sn68 3183.098862
Rwneg124_69 in124 sn69 3183.098862
Rwneg124_70 in124 sn70 3183.098862
Rwneg124_71 in124 sn71 3183.098862
Rwneg124_72 in124 sn72 3183.098862
Rwneg124_73 in124 sn73 11140.846016
Rwneg124_74 in124 sn74 11140.846016
Rwneg124_75 in124 sn75 3183.098862
Rwneg124_76 in124 sn76 3183.098862
Rwneg124_77 in124 sn77 3183.098862
Rwneg124_78 in124 sn78 3183.098862
Rwneg124_79 in124 sn79 3183.098862
Rwneg124_80 in124 sn80 11140.846016
Rwneg124_81 in124 sn81 3183.098862
Rwneg124_82 in124 sn82 3183.098862
Rwneg124_83 in124 sn83 11140.846016
Rwneg124_84 in124 sn84 11140.846016
Rwneg124_85 in124 sn85 3183.098862
Rwneg124_86 in124 sn86 3183.098862
Rwneg124_87 in124 sn87 3183.098862
Rwneg124_88 in124 sn88 11140.846016
Rwneg124_89 in124 sn89 11140.846016
Rwneg124_90 in124 sn90 3183.098862
Rwneg124_91 in124 sn91 3183.098862
Rwneg124_92 in124 sn92 3183.098862
Rwneg124_93 in124 sn93 3183.098862
Rwneg124_94 in124 sn94 11140.846016
Rwneg124_95 in124 sn95 3183.098862
Rwneg124_96 in124 sn96 3183.098862
Rwneg124_97 in124 sn97 11140.846016
Rwneg124_98 in124 sn98 3183.098862
Rwneg124_99 in124 sn99 3183.098862
Rwneg124_100 in124 sn100 11140.846016
Rwneg125_1 in125 sn1 3183.098862
Rwneg125_2 in125 sn2 11140.846016
Rwneg125_3 in125 sn3 3183.098862
Rwneg125_4 in125 sn4 3183.098862
Rwneg125_5 in125 sn5 11140.846016
Rwneg125_6 in125 sn6 3183.098862
Rwneg125_7 in125 sn7 11140.846016
Rwneg125_8 in125 sn8 11140.846016
Rwneg125_9 in125 sn9 11140.846016
Rwneg125_10 in125 sn10 11140.846016
Rwneg125_11 in125 sn11 3183.098862
Rwneg125_12 in125 sn12 11140.846016
Rwneg125_13 in125 sn13 3183.098862
Rwneg125_14 in125 sn14 11140.846016
Rwneg125_15 in125 sn15 11140.846016
Rwneg125_16 in125 sn16 3183.098862
Rwneg125_17 in125 sn17 3183.098862
Rwneg125_18 in125 sn18 3183.098862
Rwneg125_19 in125 sn19 11140.846016
Rwneg125_20 in125 sn20 11140.846016
Rwneg125_21 in125 sn21 11140.846016
Rwneg125_22 in125 sn22 3183.098862
Rwneg125_23 in125 sn23 3183.098862
Rwneg125_24 in125 sn24 11140.846016
Rwneg125_25 in125 sn25 3183.098862
Rwneg125_26 in125 sn26 3183.098862
Rwneg125_27 in125 sn27 11140.846016
Rwneg125_28 in125 sn28 11140.846016
Rwneg125_29 in125 sn29 3183.098862
Rwneg125_30 in125 sn30 3183.098862
Rwneg125_31 in125 sn31 3183.098862
Rwneg125_32 in125 sn32 3183.098862
Rwneg125_33 in125 sn33 3183.098862
Rwneg125_34 in125 sn34 3183.098862
Rwneg125_35 in125 sn35 3183.098862
Rwneg125_36 in125 sn36 11140.846016
Rwneg125_37 in125 sn37 3183.098862
Rwneg125_38 in125 sn38 11140.846016
Rwneg125_39 in125 sn39 3183.098862
Rwneg125_40 in125 sn40 11140.846016
Rwneg125_41 in125 sn41 3183.098862
Rwneg125_42 in125 sn42 3183.098862
Rwneg125_43 in125 sn43 11140.846016
Rwneg125_44 in125 sn44 3183.098862
Rwneg125_45 in125 sn45 3183.098862
Rwneg125_46 in125 sn46 3183.098862
Rwneg125_47 in125 sn47 3183.098862
Rwneg125_48 in125 sn48 3183.098862
Rwneg125_49 in125 sn49 3183.098862
Rwneg125_50 in125 sn50 11140.846016
Rwneg125_51 in125 sn51 3183.098862
Rwneg125_52 in125 sn52 3183.098862
Rwneg125_53 in125 sn53 3183.098862
Rwneg125_54 in125 sn54 11140.846016
Rwneg125_55 in125 sn55 11140.846016
Rwneg125_56 in125 sn56 11140.846016
Rwneg125_57 in125 sn57 11140.846016
Rwneg125_58 in125 sn58 3183.098862
Rwneg125_59 in125 sn59 11140.846016
Rwneg125_60 in125 sn60 3183.098862
Rwneg125_61 in125 sn61 11140.846016
Rwneg125_62 in125 sn62 11140.846016
Rwneg125_63 in125 sn63 3183.098862
Rwneg125_64 in125 sn64 11140.846016
Rwneg125_65 in125 sn65 11140.846016
Rwneg125_66 in125 sn66 3183.098862
Rwneg125_67 in125 sn67 3183.098862
Rwneg125_68 in125 sn68 3183.098862
Rwneg125_69 in125 sn69 3183.098862
Rwneg125_70 in125 sn70 11140.846016
Rwneg125_71 in125 sn71 11140.846016
Rwneg125_72 in125 sn72 3183.098862
Rwneg125_73 in125 sn73 3183.098862
Rwneg125_74 in125 sn74 11140.846016
Rwneg125_75 in125 sn75 3183.098862
Rwneg125_76 in125 sn76 11140.846016
Rwneg125_77 in125 sn77 11140.846016
Rwneg125_78 in125 sn78 3183.098862
Rwneg125_79 in125 sn79 3183.098862
Rwneg125_80 in125 sn80 3183.098862
Rwneg125_81 in125 sn81 11140.846016
Rwneg125_82 in125 sn82 3183.098862
Rwneg125_83 in125 sn83 3183.098862
Rwneg125_84 in125 sn84 11140.846016
Rwneg125_85 in125 sn85 11140.846016
Rwneg125_86 in125 sn86 11140.846016
Rwneg125_87 in125 sn87 3183.098862
Rwneg125_88 in125 sn88 11140.846016
Rwneg125_89 in125 sn89 3183.098862
Rwneg125_90 in125 sn90 11140.846016
Rwneg125_91 in125 sn91 11140.846016
Rwneg125_92 in125 sn92 3183.098862
Rwneg125_93 in125 sn93 3183.098862
Rwneg125_94 in125 sn94 3183.098862
Rwneg125_95 in125 sn95 11140.846016
Rwneg125_96 in125 sn96 11140.846016
Rwneg125_97 in125 sn97 11140.846016
Rwneg125_98 in125 sn98 11140.846016
Rwneg125_99 in125 sn99 11140.846016
Rwneg125_100 in125 sn100 11140.846016
Rwneg126_1 in126 sn1 11140.846016
Rwneg126_2 in126 sn2 11140.846016
Rwneg126_3 in126 sn3 11140.846016
Rwneg126_4 in126 sn4 3183.098862
Rwneg126_5 in126 sn5 11140.846016
Rwneg126_6 in126 sn6 11140.846016
Rwneg126_7 in126 sn7 11140.846016
Rwneg126_8 in126 sn8 3183.098862
Rwneg126_9 in126 sn9 11140.846016
Rwneg126_10 in126 sn10 11140.846016
Rwneg126_11 in126 sn11 3183.098862
Rwneg126_12 in126 sn12 11140.846016
Rwneg126_13 in126 sn13 3183.098862
Rwneg126_14 in126 sn14 3183.098862
Rwneg126_15 in126 sn15 3183.098862
Rwneg126_16 in126 sn16 11140.846016
Rwneg126_17 in126 sn17 11140.846016
Rwneg126_18 in126 sn18 11140.846016
Rwneg126_19 in126 sn19 11140.846016
Rwneg126_20 in126 sn20 11140.846016
Rwneg126_21 in126 sn21 11140.846016
Rwneg126_22 in126 sn22 3183.098862
Rwneg126_23 in126 sn23 11140.846016
Rwneg126_24 in126 sn24 3183.098862
Rwneg126_25 in126 sn25 11140.846016
Rwneg126_26 in126 sn26 3183.098862
Rwneg126_27 in126 sn27 3183.098862
Rwneg126_28 in126 sn28 3183.098862
Rwneg126_29 in126 sn29 11140.846016
Rwneg126_30 in126 sn30 3183.098862
Rwneg126_31 in126 sn31 11140.846016
Rwneg126_32 in126 sn32 11140.846016
Rwneg126_33 in126 sn33 3183.098862
Rwneg126_34 in126 sn34 3183.098862
Rwneg126_35 in126 sn35 3183.098862
Rwneg126_36 in126 sn36 11140.846016
Rwneg126_37 in126 sn37 3183.098862
Rwneg126_38 in126 sn38 11140.846016
Rwneg126_39 in126 sn39 3183.098862
Rwneg126_40 in126 sn40 11140.846016
Rwneg126_41 in126 sn41 3183.098862
Rwneg126_42 in126 sn42 11140.846016
Rwneg126_43 in126 sn43 3183.098862
Rwneg126_44 in126 sn44 11140.846016


**********Positive Biases****************

Rbpos1 vdd sp1 3183.098862
Rbpos2 vdd sp2 3183.098862
Rbpos3 vdd sp3 3183.098862
Rbpos4 vdd sp4 11140.846016
Rbpos5 vdd sp5 3183.098862
Rbpos6 vdd sp6 3183.098862
Rbpos7 vdd sp7 11140.846016
Rbpos8 vdd sp8 3183.098862
Rbpos9 vdd sp9 11140.846016
Rbpos10 vdd sp10 3183.098862
Rbpos11 vdd sp11 3183.098862
Rbpos12 vdd sp12 3183.098862
Rbpos13 vdd sp13 3183.098862
Rbpos14 vdd sp14 3183.098862
Rbpos15 vdd sp15 3183.098862
Rbpos16 vdd sp16 3183.098862


**********Negative Biases****************

Rbneg1 vss sn1 11140.846016
Rbneg2 vss sn2 11140.846016
Rbneg3 vss sn3 11140.846016
Rbneg4 vss sn4 3183.098862
Rbneg5 vss sn5 11140.846016
Rbneg6 vss sn6 11140.846016
Rbneg7 vss sn7 3183.098862
Rbneg8 vss sn8 11140.846016
Rbneg9 vss sn9 3183.098862
Rbneg10 vss sn10 11140.846016
Rbneg11 vss sn11 11140.846016
Rbneg12 vss sn12 11140.846016
Rbneg13 vss sn13 11140.846016
Rbneg14 vss sn14 11140.846016
Rbneg15 vss sn15 11140.846016
Rbneg16 vss sn16 11140.846016


**********Weight Differntial Op-AMPS****************

XDIFFw1 sp1 sn1 xin1 diff
XDIFFw2 sp2 sn2 xin2 diff
XDIFFw3 sp3 sn3 xin3 diff
XDIFFw4 sp4 sn4 xin4 diff
XDIFFw5 sp5 sn5 xin5 diff
XDIFFw6 sp6 sn6 xin6 diff
XDIFFw7 sp7 sn7 xin7 diff
XDIFFw8 sp8 sn8 xin8 diff
XDIFFw9 sp9 sn9 xin9 diff
XDIFFw10 sp10 sn10 xin10 diff
XDIFFw11 sp11 sn11 xin11 diff
XDIFFw12 sp12 sn12 xin12 diff
XDIFFw13 sp13 sn13 xin13 diff
XDIFFw14 sp14 sn14 xin14 diff
XDIFFw15 sp15 sn15 xin15 diff
XDIFFw16 sp16 sn16 xin16 diff
XDIFFw17 sp17 sn17 xin17 diff
XDIFFw18 sp18 sn18 xin18 diff
XDIFFw19 sp19 sn19 xin19 diff
XDIFFw20 sp20 sn20 xin20 diff
XDIFFw21 sp21 sn21 xin21 diff
XDIFFw22 sp22 sn22 xin22 diff
XDIFFw23 sp23 sn23 xin23 diff
XDIFFw24 sp24 sn24 xin24 diff
XDIFFw25 sp25 sn25 xin25 diff
XDIFFw26 sp26 sn26 xin26 diff
XDIFFw27 sp27 sn27 xin27 diff
XDIFFw28 sp28 sn28 xin28 diff
XDIFFw29 sp29 sn29 xin29 diff
XDIFFw30 sp30 sn30 xin30 diff
XDIFFw31 sp31 sn31 xin31 diff
XDIFFw32 sp32 sn32 xin32 diff
XDIFFw33 sp33 sn33 xin33 diff
XDIFFw34 sp34 sn34 xin34 diff
XDIFFw35 sp35 sn35 xin35 diff
XDIFFw36 sp36 sn36 xin36 diff
XDIFFw37 sp37 sn37 xin37 diff
XDIFFw38 sp38 sn38 xin38 diff
XDIFFw39 sp39 sn39 xin39 diff
XDIFFw40 sp40 sn40 xin40 diff
XDIFFw41 sp41 sn41 xin41 diff
XDIFFw42 sp42 sn42 xin42 diff
XDIFFw43 sp43 sn43 xin43 diff
XDIFFw44 sp44 sn44 xin44 diff
XDIFFw45 sp45 sn45 xin45 diff
XDIFFw46 sp46 sn46 xin46 diff
XDIFFw47 sp47 sn47 xin47 diff
XDIFFw48 sp48 sn48 xin48 diff
XDIFFw49 sp49 sn49 xin49 diff
XDIFFw50 sp50 sn50 xin50 diff
XDIFFw51 sp51 sn51 xin51 diff
XDIFFw52 sp52 sn52 xin52 diff
XDIFFw53 sp53 sn53 xin53 diff
XDIFFw54 sp54 sn54 xin54 diff
XDIFFw55 sp55 sn55 xin55 diff
XDIFFw56 sp56 sn56 xin56 diff
XDIFFw57 sp57 sn57 xin57 diff
XDIFFw58 sp58 sn58 xin58 diff
XDIFFw59 sp59 sn59 xin59 diff
XDIFFw60 sp60 sn60 xin60 diff
XDIFFw61 sp61 sn61 xin61 diff
XDIFFw62 sp62 sn62 xin62 diff
XDIFFw63 sp63 sn63 xin63 diff
XDIFFw64 sp64 sn64 xin64 diff
XDIFFw65 sp65 sn65 xin65 diff
XDIFFw66 sp66 sn66 xin66 diff
XDIFFw67 sp67 sn67 xin67 diff
XDIFFw68 sp68 sn68 xin68 diff
XDIFFw69 sp69 sn69 xin69 diff
XDIFFw70 sp70 sn70 xin70 diff
XDIFFw71 sp71 sn71 xin71 diff
XDIFFw72 sp72 sn72 xin72 diff
XDIFFw73 sp73 sn73 xin73 diff
XDIFFw74 sp74 sn74 xin74 diff
XDIFFw75 sp75 sn75 xin75 diff
XDIFFw76 sp76 sn76 xin76 diff
XDIFFw77 sp77 sn77 xin77 diff
XDIFFw78 sp78 sn78 xin78 diff
XDIFFw79 sp79 sn79 xin79 diff
XDIFFw80 sp80 sn80 xin80 diff
XDIFFw81 sp81 sn81 xin81 diff
XDIFFw82 sp82 sn82 xin82 diff
XDIFFw83 sp83 sn83 xin83 diff
XDIFFw84 sp84 sn84 xin84 diff
XDIFFw85 sp85 sn85 xin85 diff
XDIFFw86 sp86 sn86 xin86 diff
XDIFFw87 sp87 sn87 xin87 diff
XDIFFw88 sp88 sn88 xin88 diff
XDIFFw89 sp89 sn89 xin89 diff
XDIFFw90 sp90 sn90 xin90 diff
XDIFFw91 sp91 sn91 xin91 diff
XDIFFw92 sp92 sn92 xin92 diff
XDIFFw93 sp93 sn93 xin93 diff
XDIFFw94 sp94 sn94 xin94 diff
XDIFFw95 sp95 sn95 xin95 diff
XDIFFw96 sp96 sn96 xin96 diff
XDIFFw97 sp97 sn97 xin97 diff
XDIFFw98 sp98 sn98 xin98 diff
XDIFFw99 sp99 sn99 xin99 diff
XDIFFw100 sp100 sn100 xin100 diff


**********neurons****************

Xsig1 xin1 out1 vdd 0 neuron
Xsig2 xin2 out2 vdd 0 neuron
Xsig3 xin3 out3 vdd 0 neuron
Xsig4 xin4 out4 vdd 0 neuron
Xsig5 xin5 out5 vdd 0 neuron
Xsig6 xin6 out6 vdd 0 neuron
Xsig7 xin7 out7 vdd 0 neuron
Xsig8 xin8 out8 vdd 0 neuron
Xsig9 xin9 out9 vdd 0 neuron
Xsig10 xin10 out10 vdd 0 neuron
Xsig11 xin11 out11 vdd 0 neuron
Xsig12 xin12 out12 vdd 0 neuron
Xsig13 xin13 out13 vdd 0 neuron
Xsig14 xin14 out14 vdd 0 neuron
Xsig15 xin15 out15 vdd 0 neuron
Xsig16 xin16 out16 vdd 0 neuron
Xsig17 xin17 out17 vdd 0 neuron
Xsig18 xin18 out18 vdd 0 neuron
Xsig19 xin19 out19 vdd 0 neuron
Xsig20 xin20 out20 vdd 0 neuron
Xsig21 xin21 out21 vdd 0 neuron
Xsig22 xin22 out22 vdd 0 neuron
Xsig23 xin23 out23 vdd 0 neuron
Xsig24 xin24 out24 vdd 0 neuron
Xsig25 xin25 out25 vdd 0 neuron
Xsig26 xin26 out26 vdd 0 neuron
Xsig27 xin27 out27 vdd 0 neuron
Xsig28 xin28 out28 vdd 0 neuron
Xsig29 xin29 out29 vdd 0 neuron
Xsig30 xin30 out30 vdd 0 neuron
Xsig31 xin31 out31 vdd 0 neuron
Xsig32 xin32 out32 vdd 0 neuron
Xsig33 xin33 out33 vdd 0 neuron
Xsig34 xin34 out34 vdd 0 neuron
Xsig35 xin35 out35 vdd 0 neuron
Xsig36 xin36 out36 vdd 0 neuron
Xsig37 xin37 out37 vdd 0 neuron
Xsig38 xin38 out38 vdd 0 neuron
Xsig39 xin39 out39 vdd 0 neuron
Xsig40 xin40 out40 vdd 0 neuron
Xsig41 xin41 out41 vdd 0 neuron
Xsig42 xin42 out42 vdd 0 neuron
Xsig43 xin43 out43 vdd 0 neuron
Xsig44 xin44 out44 vdd 0 neuron
Xsig45 xin45 out45 vdd 0 neuron
Xsig46 xin46 out46 vdd 0 neuron
Xsig47 xin47 out47 vdd 0 neuron
Xsig48 xin48 out48 vdd 0 neuron
Xsig49 xin49 out49 vdd 0 neuron
Xsig50 xin50 out50 vdd 0 neuron
Xsig51 xin51 out51 vdd 0 neuron
Xsig52 xin52 out52 vdd 0 neuron
Xsig53 xin53 out53 vdd 0 neuron
Xsig54 xin54 out54 vdd 0 neuron
Xsig55 xin55 out55 vdd 0 neuron
Xsig56 xin56 out56 vdd 0 neuron
Xsig57 xin57 out57 vdd 0 neuron
Xsig58 xin58 out58 vdd 0 neuron
Xsig59 xin59 out59 vdd 0 neuron
Xsig60 xin60 out60 vdd 0 neuron
Xsig61 xin61 out61 vdd 0 neuron
Xsig62 xin62 out62 vdd 0 neuron
Xsig63 xin63 out63 vdd 0 neuron
Xsig64 xin64 out64 vdd 0 neuron
Xsig65 xin65 out65 vdd 0 neuron
Xsig66 xin66 out66 vdd 0 neuron
Xsig67 xin67 out67 vdd 0 neuron
Xsig68 xin68 out68 vdd 0 neuron
Xsig69 xin69 out69 vdd 0 neuron
Xsig70 xin70 out70 vdd 0 neuron
Xsig71 xin71 out71 vdd 0 neuron
Xsig72 xin72 out72 vdd 0 neuron
Xsig73 xin73 out73 vdd 0 neuron
Xsig74 xin74 out74 vdd 0 neuron
Xsig75 xin75 out75 vdd 0 neuron
Xsig76 xin76 out76 vdd 0 neuron
Xsig77 xin77 out77 vdd 0 neuron
Xsig78 xin78 out78 vdd 0 neuron
Xsig79 xin79 out79 vdd 0 neuron
Xsig80 xin80 out80 vdd 0 neuron
Xsig81 xin81 out81 vdd 0 neuron
Xsig82 xin82 out82 vdd 0 neuron
Xsig83 xin83 out83 vdd 0 neuron
Xsig84 xin84 out84 vdd 0 neuron
Xsig85 xin85 out85 vdd 0 neuron
Xsig86 xin86 out86 vdd 0 neuron
Xsig87 xin87 out87 vdd 0 neuron
Xsig88 xin88 out88 vdd 0 neuron
Xsig89 xin89 out89 vdd 0 neuron
Xsig90 xin90 out90 vdd 0 neuron
Xsig91 xin91 out91 vdd 0 neuron
Xsig92 xin92 out92 vdd 0 neuron
Xsig93 xin93 out93 vdd 0 neuron
Xsig94 xin94 out94 vdd 0 neuron
Xsig95 xin95 out95 vdd 0 neuron
Xsig96 xin96 out96 vdd 0 neuron
Xsig97 xin97 out97 vdd 0 neuron
Xsig98 xin98 out98 vdd 0 neuron
Xsig99 xin99 out99 vdd 0 neuron
Xsig100 xin100 out100 vdd 0 neuron
.ENDS layer1
.SUBCKT layer2 vdd vss in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15 in16 in17 in18 in19 in20 in21 in22 in23 in24 in25 in26 in27 in28 in29 in30 in31 in32 in33 in34 in35 in36 in37 in38 in39 in40 in41 in42 in43 in44 in45 in46 in47 in48 in49 in50 in51 in52 in53 in54 in55 in56 in57 in58 in59 in60 in61 in62 in63 in64 in65 in66 in67 in68 in69 in70 in71 in72 in73 in74 in75 in76 in77 in78 in79 in80 in81 in82 in83 in84 in85 in86 in87 in88 in89 in90 in91 in92 in93 in94 in95 in96 in97 in98 in99 in100 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 

**********Non-Negative Weighted Array****************
Rwpos1_1 in1 sp1 3183.098862
Rwpos1_2 in1 sp2 3183.098862
Rwpos1_3 in1 sp3 3183.098862
Rwpos1_4 in1 sp4 11140.846016
Rwpos1_5 in1 sp5 3183.098862
Rwpos1_6 in1 sp6 3183.098862
Rwpos1_7 in1 sp7 3183.098862
Rwpos1_8 in1 sp8 11140.846016
Rwpos1_9 in1 sp9 3183.098862
Rwpos1_10 in1 sp10 3183.098862
Rwpos2_1 in2 sp1 3183.098862
Rwpos2_2 in2 sp2 3183.098862
Rwpos2_3 in2 sp3 3183.098862
Rwpos2_4 in2 sp4 11140.846016
Rwpos2_5 in2 sp5 11140.846016
Rwpos2_6 in2 sp6 3183.098862
Rwpos2_7 in2 sp7 3183.098862
Rwpos2_8 in2 sp8 3183.098862
Rwpos2_9 in2 sp9 11140.846016
Rwpos2_10 in2 sp10 3183.098862
Rwpos3_1 in3 sp1 3183.098862
Rwpos3_2 in3 sp2 3183.098862
Rwpos3_3 in3 sp3 3183.098862
Rwpos3_4 in3 sp4 3183.098862
Rwpos3_5 in3 sp5 3183.098862
Rwpos3_6 in3 sp6 3183.098862
Rwpos3_7 in3 sp7 3183.098862
Rwpos3_8 in3 sp8 3183.098862
Rwpos3_9 in3 sp9 3183.098862
Rwpos3_10 in3 sp10 11140.846016
Rwpos4_1 in4 sp1 3183.098862
Rwpos4_2 in4 sp2 11140.846016
Rwpos4_3 in4 sp3 3183.098862
Rwpos4_4 in4 sp4 3183.098862
Rwpos4_5 in4 sp5 3183.098862
Rwpos4_6 in4 sp6 3183.098862
Rwpos4_7 in4 sp7 3183.098862
Rwpos4_8 in4 sp8 11140.846016
Rwpos4_9 in4 sp9 3183.098862
Rwpos4_10 in4 sp10 3183.098862
Rwpos5_1 in5 sp1 3183.098862
Rwpos5_2 in5 sp2 3183.098862
Rwpos5_3 in5 sp3 11140.846016
Rwpos5_4 in5 sp4 3183.098862
Rwpos5_5 in5 sp5 3183.098862
Rwpos5_6 in5 sp6 3183.098862
Rwpos5_7 in5 sp7 3183.098862
Rwpos5_8 in5 sp8 11140.846016
Rwpos5_9 in5 sp9 3183.098862
Rwpos5_10 in5 sp10 3183.098862
Rwpos6_1 in6 sp1 3183.098862
Rwpos6_2 in6 sp2 3183.098862
Rwpos6_3 in6 sp3 3183.098862
Rwpos6_4 in6 sp4 11140.846016
Rwpos6_5 in6 sp5 3183.098862
Rwpos6_6 in6 sp6 3183.098862
Rwpos6_7 in6 sp7 11140.846016
Rwpos6_8 in6 sp8 3183.098862
Rwpos6_9 in6 sp9 3183.098862
Rwpos6_10 in6 sp10 3183.098862
Rwpos7_1 in7 sp1 3183.098862
Rwpos7_2 in7 sp2 11140.846016
Rwpos7_3 in7 sp3 3183.098862
Rwpos7_4 in7 sp4 3183.098862
Rwpos7_5 in7 sp5 3183.098862
Rwpos7_6 in7 sp6 11140.846016
Rwpos7_7 in7 sp7 3183.098862
Rwpos7_8 in7 sp8 3183.098862
Rwpos7_9 in7 sp9 3183.098862
Rwpos7_10 in7 sp10 3183.098862
Rwpos8_1 in8 sp1 3183.098862
Rwpos8_2 in8 sp2 3183.098862
Rwpos8_3 in8 sp3 3183.098862
Rwpos8_4 in8 sp4 3183.098862
Rwpos8_5 in8 sp5 11140.846016
Rwpos8_6 in8 sp6 3183.098862
Rwpos8_7 in8 sp7 3183.098862
Rwpos8_8 in8 sp8 3183.098862
Rwpos8_9 in8 sp9 3183.098862
Rwpos8_10 in8 sp10 11140.846016
Rwpos9_1 in9 sp1 11140.846016
Rwpos9_2 in9 sp2 3183.098862
Rwpos9_3 in9 sp3 3183.098862
Rwpos9_4 in9 sp4 3183.098862
Rwpos9_5 in9 sp5 3183.098862
Rwpos9_6 in9 sp6 11140.846016
Rwpos9_7 in9 sp7 11140.846016
Rwpos9_8 in9 sp8 3183.098862
Rwpos9_9 in9 sp9 3183.098862
Rwpos9_10 in9 sp10 3183.098862
Rwpos10_1 in10 sp1 3183.098862
Rwpos10_2 in10 sp2 3183.098862
Rwpos10_3 in10 sp3 3183.098862
Rwpos10_4 in10 sp4 3183.098862
Rwpos10_5 in10 sp5 11140.846016
Rwpos10_6 in10 sp6 3183.098862
Rwpos10_7 in10 sp7 11140.846016
Rwpos10_8 in10 sp8 3183.098862
Rwpos10_9 in10 sp9 3183.098862
Rwpos10_10 in10 sp10 3183.098862
Rwpos11_1 in11 sp1 3183.098862
Rwpos11_2 in11 sp2 3183.098862
Rwpos11_3 in11 sp3 11140.846016
Rwpos11_4 in11 sp4 11140.846016
Rwpos11_5 in11 sp5 3183.098862
Rwpos11_6 in11 sp6 3183.098862
Rwpos11_7 in11 sp7 3183.098862
Rwpos11_8 in11 sp8 3183.098862
Rwpos11_9 in11 sp9 3183.098862
Rwpos11_10 in11 sp10 3183.098862
Rwpos12_1 in12 sp1 11140.846016
Rwpos12_2 in12 sp2 3183.098862
Rwpos12_3 in12 sp3 11140.846016
Rwpos12_4 in12 sp4 3183.098862
Rwpos12_5 in12 sp5 3183.098862
Rwpos12_6 in12 sp6 3183.098862
Rwpos12_7 in12 sp7 3183.098862
Rwpos12_8 in12 sp8 3183.098862
Rwpos12_9 in12 sp9 3183.098862
Rwpos12_10 in12 sp10 3183.098862
Rwpos13_1 in13 sp1 3183.098862
Rwpos13_2 in13 sp2 3183.098862
Rwpos13_3 in13 sp3 3183.098862
Rwpos13_4 in13 sp4 3183.098862
Rwpos13_5 in13 sp5 3183.098862
Rwpos13_6 in13 sp6 11140.846016
Rwpos13_7 in13 sp7 3183.098862
Rwpos13_8 in13 sp8 3183.098862
Rwpos13_9 in13 sp9 11140.846016
Rwpos13_10 in13 sp10 3183.098862
Rwpos14_1 in14 sp1 3183.098862
Rwpos14_2 in14 sp2 11140.846016
Rwpos14_3 in14 sp3 11140.846016
Rwpos14_4 in14 sp4 3183.098862
Rwpos14_5 in14 sp5 3183.098862
Rwpos14_6 in14 sp6 3183.098862
Rwpos14_7 in14 sp7 3183.098862
Rwpos14_8 in14 sp8 3183.098862
Rwpos14_9 in14 sp9 11140.846016
Rwpos14_10 in14 sp10 3183.098862
Rwpos15_1 in15 sp1 11140.846016
Rwpos15_2 in15 sp2 3183.098862
Rwpos15_3 in15 sp3 3183.098862
Rwpos15_4 in15 sp4 3183.098862
Rwpos15_5 in15 sp5 3183.098862
Rwpos15_6 in15 sp6 3183.098862
Rwpos15_7 in15 sp7 3183.098862
Rwpos15_8 in15 sp8 11140.846016
Rwpos15_9 in15 sp9 3183.098862
Rwpos15_10 in15 sp10 3183.098862
Rwpos16_1 in16 sp1 3183.098862
Rwpos16_2 in16 sp2 3183.098862
Rwpos16_3 in16 sp3 11140.846016
Rwpos16_4 in16 sp4 3183.098862
Rwpos16_5 in16 sp5 3183.098862
Rwpos16_6 in16 sp6 3183.098862
Rwpos16_7 in16 sp7 11140.846016
Rwpos16_8 in16 sp8 3183.098862
Rwpos16_9 in16 sp9 3183.098862
Rwpos16_10 in16 sp10 3183.098862


**********Negative Weighted Array****************

Rwneg1_1 in1 sn1 11140.846016
Rwneg1_2 in1 sn2 11140.846016
Rwneg1_3 in1 sn3 11140.846016
Rwneg1_4 in1 sn4 3183.098862
Rwneg1_5 in1 sn5 11140.846016
Rwneg1_6 in1 sn6 11140.846016
Rwneg1_7 in1 sn7 11140.846016
Rwneg1_8 in1 sn8 3183.098862
Rwneg1_9 in1 sn9 11140.846016
Rwneg1_10 in1 sn10 11140.846016
Rwneg2_1 in2 sn1 11140.846016
Rwneg2_2 in2 sn2 11140.846016
Rwneg2_3 in2 sn3 11140.846016
Rwneg2_4 in2 sn4 3183.098862
Rwneg2_5 in2 sn5 3183.098862
Rwneg2_6 in2 sn6 11140.846016
Rwneg2_7 in2 sn7 11140.846016
Rwneg2_8 in2 sn8 11140.846016
Rwneg2_9 in2 sn9 3183.098862
Rwneg2_10 in2 sn10 11140.846016
Rwneg3_1 in3 sn1 11140.846016
Rwneg3_2 in3 sn2 11140.846016
Rwneg3_3 in3 sn3 11140.846016
Rwneg3_4 in3 sn4 11140.846016
Rwneg3_5 in3 sn5 11140.846016
Rwneg3_6 in3 sn6 11140.846016
Rwneg3_7 in3 sn7 11140.846016
Rwneg3_8 in3 sn8 11140.846016
Rwneg3_9 in3 sn9 11140.846016
Rwneg3_10 in3 sn10 3183.098862
Rwneg4_1 in4 sn1 11140.846016
Rwneg4_2 in4 sn2 3183.098862
Rwneg4_3 in4 sn3 11140.846016
Rwneg4_4 in4 sn4 11140.846016
Rwneg4_5 in4 sn5 11140.846016
Rwneg4_6 in4 sn6 11140.846016
Rwneg4_7 in4 sn7 11140.846016
Rwneg4_8 in4 sn8 3183.098862
Rwneg4_9 in4 sn9 11140.846016
Rwneg4_10 in4 sn10 11140.846016
Rwneg5_1 in5 sn1 11140.846016
Rwneg5_2 in5 sn2 11140.846016
Rwneg5_3 in5 sn3 3183.098862
Rwneg5_4 in5 sn4 11140.846016
Rwneg5_5 in5 sn5 11140.846016
Rwneg5_6 in5 sn6 11140.846016
Rwneg5_7 in5 sn7 11140.846016
Rwneg5_8 in5 sn8 3183.098862
Rwneg5_9 in5 sn9 11140.846016
Rwneg5_10 in5 sn10 11140.846016
Rwneg6_1 in6 sn1 11140.846016
Rwneg6_2 in6 sn2 11140.846016
Rwneg6_3 in6 sn3 11140.846016
Rwneg6_4 in6 sn4 3183.098862
Rwneg6_5 in6 sn5 11140.846016
Rwneg6_6 in6 sn6 11140.846016
Rwneg6_7 in6 sn7 3183.098862
Rwneg6_8 in6 sn8 11140.846016
Rwneg6_9 in6 sn9 11140.846016
Rwneg6_10 in6 sn10 11140.846016
Rwneg7_1 in7 sn1 11140.846016
Rwneg7_2 in7 sn2 3183.098862
Rwneg7_3 in7 sn3 11140.846016
Rwneg7_4 in7 sn4 11140.846016
Rwneg7_5 in7 sn5 11140.846016
Rwneg7_6 in7 sn6 3183.098862
Rwneg7_7 in7 sn7 11140.846016
Rwneg7_8 in7 sn8 11140.846016
Rwneg7_9 in7 sn9 11140.846016
Rwneg7_10 in7 sn10 11140.846016
Rwneg8_1 in8 sn1 11140.846016
Rwneg8_2 in8 sn2 11140.846016
Rwneg8_3 in8 sn3 11140.846016
Rwneg8_4 in8 sn4 11140.846016
Rwneg8_5 in8 sn5 3183.098862
Rwneg8_6 in8 sn6 11140.846016
Rwneg8_7 in8 sn7 11140.846016
Rwneg8_8 in8 sn8 11140.846016
Rwneg8_9 in8 sn9 11140.846016
Rwneg8_10 in8 sn10 3183.098862
Rwneg9_1 in9 sn1 3183.098862
Rwneg9_2 in9 sn2 11140.846016
Rwneg9_3 in9 sn3 11140.846016
Rwneg9_4 in9 sn4 11140.846016
Rwneg9_5 in9 sn5 11140.846016
Rwneg9_6 in9 sn6 3183.098862
Rwneg9_7 in9 sn7 3183.098862
Rwneg9_8 in9 sn8 11140.846016
Rwneg9_9 in9 sn9 11140.846016
Rwneg9_10 in9 sn10 11140.846016
Rwneg10_1 in10 sn1 11140.846016
Rwneg10_2 in10 sn2 11140.846016
Rwneg10_3 in10 sn3 11140.846016
Rwneg10_4 in10 sn4 11140.846016
Rwneg10_5 in10 sn5 3183.098862
Rwneg10_6 in10 sn6 11140.846016
Rwneg10_7 in10 sn7 3183.098862
Rwneg10_8 in10 sn8 11140.846016
Rwneg10_9 in10 sn9 11140.846016
Rwneg10_10 in10 sn10 11140.846016
Rwneg11_1 in11 sn1 11140.846016
Rwneg11_2 in11 sn2 11140.846016
Rwneg11_3 in11 sn3 3183.098862
Rwneg11_4 in11 sn4 3183.098862
Rwneg11_5 in11 sn5 11140.846016
Rwneg11_6 in11 sn6 11140.846016
Rwneg11_7 in11 sn7 11140.846016
Rwneg11_8 in11 sn8 11140.846016
Rwneg11_9 in11 sn9 11140.846016
Rwneg11_10 in11 sn10 11140.846016
Rwneg12_1 in12 sn1 3183.098862
Rwneg12_2 in12 sn2 11140.846016
Rwneg12_3 in12 sn3 3183.098862
Rwneg12_4 in12 sn4 11140.846016
Rwneg12_5 in12 sn5 11140.846016
Rwneg12_6 in12 sn6 11140.846016
Rwneg12_7 in12 sn7 11140.846016
Rwneg12_8 in12 sn8 11140.846016
Rwneg12_9 in12 sn9 11140.846016
Rwneg12_10 in12 sn10 11140.846016
Rwneg13_1 in13 sn1 11140.846016
Rwneg13_2 in13 sn2 11140.846016
Rwneg13_3 in13 sn3 11140.846016
Rwneg13_4 in13 sn4 11140.846016
Rwneg13_5 in13 sn5 11140.846016
Rwneg13_6 in13 sn6 3183.098862
Rwneg13_7 in13 sn7 11140.846016
Rwneg13_8 in13 sn8 11140.846016
Rwneg13_9 in13 sn9 3183.098862
Rwneg13_10 in13 sn10 11140.846016
Rwneg14_1 in14 sn1 11140.846016
Rwneg14_2 in14 sn2 3183.098862
Rwneg14_3 in14 sn3 3183.098862
Rwneg14_4 in14 sn4 11140.846016
Rwneg14_5 in14 sn5 11140.846016
Rwneg14_6 in14 sn6 11140.846016
Rwneg14_7 in14 sn7 11140.846016
Rwneg14_8 in14 sn8 11140.846016
Rwneg14_9 in14 sn9 3183.098862
Rwneg14_10 in14 sn10 11140.846016
Rwneg15_1 in15 sn1 3183.098862
Rwneg15_2 in15 sn2 11140.846016
Rwneg15_3 in15 sn3 11140.846016
Rwneg15_4 in15 sn4 11140.846016
Rwneg15_5 in15 sn5 11140.846016
Rwneg15_6 in15 sn6 11140.846016
Rwneg15_7 in15 sn7 11140.846016
Rwneg15_8 in15 sn8 3183.098862
Rwneg15_9 in15 sn9 11140.846016
Rwneg15_10 in15 sn10 11140.846016
Rwneg16_1 in16 sn1 11140.846016
Rwneg16_2 in16 sn2 11140.846016
Rwneg16_3 in16 sn3 3183.098862
Rwneg16_4 in16 sn4 11140.846016
Rwneg16_5 in16 sn5 11140.846016
Rwneg16_6 in16 sn6 11140.846016
Rwneg16_7 in16 sn7 3183.098862
Rwneg16_8 in16 sn8 11140.846016
Rwneg16_9 in16 sn9 11140.846016
Rwneg16_10 in16 sn10 11140.846016


**********Positive Biases****************

Rbpos1 vdd sp1 3183.098862
Rbpos2 vdd sp2 3183.098862
Rbpos3 vdd sp3 3183.098862
Rbpos4 vdd sp4 3183.098862
Rbpos5 vdd sp5 3183.098862
Rbpos6 vdd sp6 3183.098862
Rbpos7 vdd sp7 3183.098862
Rbpos8 vdd sp8 3183.098862
Rbpos9 vdd sp9 3183.098862
Rbpos10 vdd sp10 3183.098862


**********Negative Biases****************

Rbneg1 vss sn1 11140.846016
Rbneg2 vss sn2 11140.846016
Rbneg3 vss sn3 11140.846016
Rbneg4 vss sn4 11140.846016
Rbneg5 vss sn5 11140.846016
Rbneg6 vss sn6 11140.846016
Rbneg7 vss sn7 11140.846016
Rbneg8 vss sn8 11140.846016
Rbneg9 vss sn9 11140.846016
Rbneg10 vss sn10 11140.846016


**********Weight Differntial Op-AMPS****************

XDIFFw1 sp1 sn1 xin1 diff2
XDIFFw2 sp2 sn2 xin2 diff2
XDIFFw3 sp3 sn3 xin3 diff2
XDIFFw4 sp4 sn4 xin4 diff2
XDIFFw5 sp5 sn5 xin5 diff2
XDIFFw6 sp6 sn6 xin6 diff2
XDIFFw7 sp7 sn7 xin7 diff2
XDIFFw8 sp8 sn8 xin8 diff2
XDIFFw9 sp9 sn9 xin9 diff2
XDIFFw10 sp10 sn10 xin10 diff2


**********neurons****************

Xsig1 xin1 out1 vdd 0 neuron
Xsig2 xin2 out2 vdd 0 neuron
Xsig3 xin3 out3 vdd 0 neuron
Xsig4 xin4 out4 vdd 0 neuron
Xsig5 xin5 out5 vdd 0 neuron
Xsig6 xin6 out6 vdd 0 neuron
Xsig7 xin7 out7 vdd 0 neuron
Xsig8 xin8 out8 vdd 0 neuron
Xsig9 xin9 out9 vdd 0 neuron
Xsig10 xin10 out10 vdd 0 neuron
.ENDS layer2
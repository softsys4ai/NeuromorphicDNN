*Fully-connected Classifier
.lib './models' ptm14hp
.include 'diff.sp'
.include 'diff2.sp'
.include 'neuron.sp'
.option post
.op
.PARAM VddVal=0.8
.PARAM VssVal=-0.8
.PARAM tsampling=1n
.include 'layer1.sp'
.include 'layer2.sp'
Xlayer1 vdd vss in0 in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15 in16 in17 in18 in19 in20 in21 in22 in23 in24 in25 in26 in27 in28 in29 in30 in31 in32 in33 in34 in35 in36 in37 in38 in39 in40 in41 in42 in43 in44 in45 in46 in47 in48 in49 in50 in51 in52 in53 in54 in55 in56 in57 in58 in59 in60 in61 in62 in63 in64 in65 in66 in67 in68 in69 in70 in71 in72 in73 in74 in75 in76 in77 in78 in79 in80 in81 in82 in83 in84 in85 in86 in87 in88 in89 in90 in91 in92 in93 in94 in95 in96 in97 in98 in99 in100 in101 in102 in103 in104 in105 in106 in107 in108 in109 in110 in111 in112 in113 in114 in115 in116 in117 in118 in119 in120 in121 in122 in123 in124 in125 in126 in127 in128 in129 in130 in131 in132 in133 in134 in135 in136 in137 in138 in139 in140 in141 in142 in143 in144 in145 in146 in147 in148 in149 in150 in151 in152 in153 in154 in155 in156 in157 in158 in159 in160 in161 in162 in163 in164 in165 in166 in167 in168 in169 in170 in171 in172 in173 in174 in175 in176 in177 in178 in179 in180 in181 in182 in183 in184 in185 in186 in187 in188 in189 in190 in191 in192 in193 in194 in195 in196 in197 in198 in199 in200 in201 in202 in203 in204 in205 in206 in207 in208 in209 in210 in211 in212 in213 in214 in215 in216 in217 in218 in219 in220 in221 in222 in223 in224 in225 in226 in227 in228 in229 in230 in231 in232 in233 in234 in235 in236 in237 in238 in239 in240 in241 in242 in243 in244 in245 in246 in247 in248 in249 in250 in251 in252 in253 in254 in255 in256 in257 in258 in259 in260 in261 in262 in263 in264 in265 in266 in267 in268 in269 in270 in271 in272 in273 in274 in275 in276 in277 in278 in279 in280 in281 in282 in283 in284 in285 in286 in287 in288 in289 in290 in291 in292 in293 in294 in295 in296 in297 in298 in299 in300 in301 in302 in303 in304 in305 in306 in307 in308 in309 in310 in311 in312 in313 in314 in315 in316 in317 in318 in319 in320 in321 in322 in323 in324 in325 in326 in327 in328 in329 in330 in331 in332 in333 in334 in335 in336 in337 in338 in339 in340 in341 in342 in343 in344 in345 in346 in347 in348 in349 in350 in351 in352 in353 in354 in355 in356 in357 in358 in359 in360 in361 in362 in363 in364 in365 in366 in367 in368 in369 in370 in371 in372 in373 in374 in375 in376 in377 in378 in379 in380 in381 in382 in383 in384 in385 in386 in387 in388 in389 in390 in391 in392 in393 in394 in395 in396 in397 in398 in399 in400 in401 in402 in403 in404 in405 in406 in407 in408 in409 in410 in411 in412 in413 in414 in415 in416 in417 in418 in419 in420 in421 in422 in423 in424 in425 in426 in427 in428 in429 in430 in431 in432 in433 in434 in435 in436 in437 in438 in439 in440 in441 in442 in443 in444 in445 in446 in447 in448 in449 in450 in451 in452 in453 in454 in455 in456 in457 in458 in459 in460 in461 in462 in463 in464 in465 in466 in467 in468 in469 in470 in471 in472 in473 in474 in475 in476 in477 in478 in479 in480 in481 in482 in483 in484 in485 in486 in487 in488 in489 in490 in491 in492 in493 in494 in495 in496 in497 in498 in499 in500 in501 in502 in503 in504 in505 in506 in507 in508 in509 in510 in511 in512 in513 in514 in515 in516 in517 in518 in519 in520 in521 in522 in523 in524 in525 in526 in527 in528 in529 in530 in531 in532 in533 in534 in535 in536 in537 in538 in539 in540 in541 in542 in543 in544 in545 in546 in547 in548 in549 in550 in551 in552 in553 in554 in555 in556 in557 in558 in559 in560 in561 in562 in563 in564 in565 in566 in567 in568 in569 in570 in571 in572 in573 in574 in575 in576 in577 in578 in579 in580 in581 in582 in583 in584 in585 in586 in587 in588 in589 in590 in591 in592 in593 in594 in595 in596 in597 in598 in599 in600 in601 in602 in603 in604 in605 in606 in607 in608 in609 in610 in611 in612 in613 in614 in615 in616 in617 in618 in619 in620 in621 in622 in623 in624 in625 in626 in627 in628 in629 in630 in631 in632 in633 in634 in635 in636 in637 in638 in639 in640 in641 in642 in643 in644 in645 in646 in647 in648 in649 in650 in651 in652 in653 in654 in655 in656 in657 in658 in659 in660 in661 in662 in663 in664 in665 in666 in667 in668 in669 in670 in671 in672 in673 in674 in675 in676 in677 in678 in679 in680 in681 in682 in683 in684 in685 in686 in687 in688 in689 in690 in691 in692 in693 in694 in695 in696 in697 in698 in699 in700 in701 in702 in703 in704 in705 in706 in707 in708 in709 in710 in711 in712 in713 in714 in715 in716 in717 in718 in719 in720 in721 in722 in723 in724 in725 in726 in727 in728 in729 in730 in731 in732 in733 in734 in735 in736 in737 in738 in739 in740 in741 in742 in743 in744 in745 in746 in747 in748 in749 in750 in751 in752 in753 in754 in755 in756 in757 in758 in759 in760 in761 in762 in763 in764 in765 in766 in767 in768 in769 in770 in771 in772 in773 in774 in775 in776 in777 in778 in779 in780 in781 in782 in783 out1_0 out1_1 out1_2 out1_3 out1_4 out1_5 out1_6 out1_7 out1_8 out1_9 out1_10 out1_11 out1_12 out1_13 out1_14 out1_15 out1_16 out1_17 out1_18 out1_19 out1_20 out1_21 out1_22 out1_23 out1_24 out1_25 out1_26 out1_27 out1_28 out1_29 out1_30 out1_31 out1_32 out1_33 out1_34 out1_35 out1_36 out1_37 out1_38 out1_39 out1_40 out1_41 out1_42 out1_43 out1_44 out1_45 out1_46 out1_47 out1_48 out1_49 out1_50 out1_51 out1_52 out1_53 out1_54 out1_55 out1_56 out1_57 out1_58 out1_59 out1_60 out1_61 out1_62 out1_63 out1_64 out1_65 out1_66 out1_67 out1_68 out1_69 out1_70 out1_71 out1_72 out1_73 out1_74 out1_75 out1_76 out1_77 out1_78 out1_79 out1_80 out1_81 out1_82 out1_83 out1_84 out1_85 out1_86 out1_87 out1_88 out1_89 out1_90 out1_91 out1_92 out1_93 out1_94 out1_95 out1_96 out1_97 out1_98 out1_99 layer1


Xlayer2 vdd vss out1_0 out1_1 out1_2 out1_3 out1_4 out1_5 out1_6 out1_7 out1_8 out1_9 out1_10 out1_11 out1_12 out1_13 out1_14 out1_15 out1_16 out1_17 out1_18 out1_19 out1_20 out1_21 out1_22 out1_23 out1_24 out1_25 out1_26 out1_27 out1_28 out1_29 out1_30 out1_31 out1_32 out1_33 out1_34 out1_35 out1_36 out1_37 out1_38 out1_39 out1_40 out1_41 out1_42 out1_43 out1_44 out1_45 out1_46 out1_47 out1_48 out1_49 out1_50 out1_51 out1_52 out1_53 out1_54 out1_55 out1_56 out1_57 out1_58 out1_59 out1_60 out1_61 out1_62 out1_63 out1_64 out1_65 out1_66 out1_67 out1_68 out1_69 out1_70 out1_71 out1_72 out1_73 out1_74 out1_75 out1_76 out1_77 out1_78 out1_79 out1_80 out1_81 out1_82 out1_83 out1_84 out1_85 out1_86 out1_87 out1_88 out1_89 out1_90 out1_91 out1_92 out1_93 out1_94 out1_95 out1_96 out1_97 out1_98 out1_99 output0 output1 output2 output3 output4 output5 output6 output7 output8 output9 layer2




**********Input Test****************

v0 in0 0 DC -0.800000
v1 in1 0 DC -0.800000
v2 in2 0 DC -0.800000
v3 in3 0 DC -0.800000
v4 in4 0 DC -0.800000
v5 in5 0 DC -0.800000
v6 in6 0 DC -0.800000
v7 in7 0 DC -0.800000
v8 in8 0 DC -0.800000
v9 in9 0 DC -0.800000
v10 in10 0 DC -0.800000
v11 in11 0 DC -0.800000
v12 in12 0 DC -0.800000
v13 in13 0 DC -0.800000
v14 in14 0 DC -0.800000
v15 in15 0 DC -0.800000
v16 in16 0 DC -0.800000
v17 in17 0 DC -0.800000
v18 in18 0 DC -0.800000
v19 in19 0 DC -0.800000
v20 in20 0 DC -0.800000
v21 in21 0 DC -0.800000
v22 in22 0 DC -0.800000
v23 in23 0 DC -0.800000
v24 in24 0 DC -0.800000
v25 in25 0 DC -0.800000
v26 in26 0 DC -0.800000
v27 in27 0 DC -0.800000
v28 in28 0 DC -0.800000
v29 in29 0 DC -0.800000
v30 in30 0 DC -0.800000
v31 in31 0 DC -0.800000
v32 in32 0 DC -0.800000
v33 in33 0 DC -0.800000
v34 in34 0 DC -0.800000
v35 in35 0 DC -0.800000
v36 in36 0 DC -0.800000
v37 in37 0 DC -0.800000
v38 in38 0 DC -0.800000
v39 in39 0 DC -0.800000
v40 in40 0 DC -0.800000
v41 in41 0 DC -0.800000
v42 in42 0 DC -0.800000
v43 in43 0 DC -0.800000
v44 in44 0 DC -0.800000
v45 in45 0 DC -0.800000
v46 in46 0 DC -0.800000
v47 in47 0 DC -0.800000
v48 in48 0 DC -0.800000
v49 in49 0 DC -0.800000
v50 in50 0 DC -0.800000
v51 in51 0 DC -0.800000
v52 in52 0 DC -0.800000
v53 in53 0 DC -0.800000
v54 in54 0 DC -0.800000
v55 in55 0 DC -0.800000
v56 in56 0 DC -0.800000
v57 in57 0 DC -0.800000
v58 in58 0 DC -0.800000
v59 in59 0 DC -0.800000
v60 in60 0 DC -0.800000
v61 in61 0 DC -0.800000
v62 in62 0 DC -0.800000
v63 in63 0 DC -0.800000
v64 in64 0 DC -0.800000
v65 in65 0 DC -0.800000
v66 in66 0 DC -0.800000
v67 in67 0 DC -0.800000
v68 in68 0 DC -0.800000
v69 in69 0 DC -0.800000
v70 in70 0 DC -0.800000
v71 in71 0 DC -0.800000
v72 in72 0 DC -0.800000
v73 in73 0 DC -0.800000
v74 in74 0 DC -0.800000
v75 in75 0 DC -0.800000
v76 in76 0 DC -0.800000
v77 in77 0 DC -0.800000
v78 in78 0 DC -0.800000
v79 in79 0 DC -0.800000
v80 in80 0 DC -0.800000
v81 in81 0 DC -0.800000
v82 in82 0 DC -0.800000
v83 in83 0 DC -0.800000
v84 in84 0 DC -0.800000
v85 in85 0 DC -0.800000
v86 in86 0 DC -0.800000
v87 in87 0 DC -0.800000
v88 in88 0 DC -0.800000
v89 in89 0 DC -0.800000
v90 in90 0 DC -0.800000
v91 in91 0 DC -0.800000
v92 in92 0 DC -0.800000
v93 in93 0 DC -0.800000
v94 in94 0 DC -0.800000
v95 in95 0 DC -0.800000
v96 in96 0 DC -0.800000
v97 in97 0 DC -0.800000
v98 in98 0 DC -0.800000
v99 in99 0 DC -0.800000
v100 in100 0 DC -0.800000
v101 in101 0 DC -0.800000
v102 in102 0 DC -0.800000
v103 in103 0 DC -0.800000
v104 in104 0 DC -0.800000
v105 in105 0 DC -0.800000
v106 in106 0 DC -0.800000
v107 in107 0 DC -0.800000
v108 in108 0 DC -0.800000
v109 in109 0 DC -0.800000
v110 in110 0 DC -0.800000
v111 in111 0 DC -0.800000
v112 in112 0 DC -0.800000
v113 in113 0 DC -0.800000
v114 in114 0 DC -0.800000
v115 in115 0 DC -0.800000
v116 in116 0 DC -0.800000
v117 in117 0 DC -0.800000
v118 in118 0 DC -0.800000
v119 in119 0 DC -0.800000
v120 in120 0 DC -0.800000
v121 in121 0 DC -0.800000
v122 in122 0 DC -0.800000
v123 in123 0 DC -0.800000
v124 in124 0 DC -0.730981
v125 in125 0 DC 0.141176
v126 in126 0 DC 0.787451
v127 in127 0 DC 0.467451
v128 in128 0 DC -0.605490
v129 in129 0 DC -0.800000
v130 in130 0 DC -0.800000
v131 in131 0 DC -0.800000
v132 in132 0 DC -0.800000
v133 in133 0 DC -0.800000
v134 in134 0 DC -0.800000
v135 in135 0 DC -0.800000
v136 in136 0 DC -0.800000
v137 in137 0 DC -0.800000
v138 in138 0 DC -0.800000
v139 in139 0 DC -0.800000
v140 in140 0 DC -0.800000
v141 in141 0 DC -0.800000
v142 in142 0 DC -0.800000
v143 in143 0 DC -0.800000
v144 in144 0 DC -0.800000
v145 in145 0 DC -0.800000
v146 in146 0 DC -0.800000
v147 in147 0 DC -0.800000
v148 in148 0 DC -0.800000
v149 in149 0 DC -0.800000
v150 in150 0 DC -0.800000
v151 in151 0 DC -0.800000
v152 in152 0 DC -0.567843
v153 in153 0 DC 0.774902
v154 in154 0 DC 0.774902
v155 in155 0 DC 0.787451
v156 in156 0 DC -0.128627
v157 in157 0 DC -0.800000
v158 in158 0 DC -0.800000
v159 in159 0 DC -0.800000
v160 in160 0 DC -0.800000
v161 in161 0 DC -0.800000
v162 in162 0 DC -0.800000
v163 in163 0 DC -0.800000
v164 in164 0 DC -0.800000
v165 in165 0 DC -0.800000
v166 in166 0 DC -0.800000
v167 in167 0 DC -0.800000
v168 in168 0 DC -0.800000
v169 in169 0 DC -0.800000
v170 in170 0 DC -0.800000
v171 in171 0 DC -0.800000
v172 in172 0 DC -0.800000
v173 in173 0 DC -0.800000
v174 in174 0 DC -0.800000
v175 in175 0 DC -0.800000
v176 in176 0 DC -0.800000
v177 in177 0 DC -0.800000
v178 in178 0 DC -0.800000
v179 in179 0 DC -0.668235
v180 in180 0 DC 0.436078
v181 in181 0 DC 0.774902
v182 in182 0 DC 0.774902
v183 in183 0 DC 0.787451
v184 in184 0 DC -0.128627
v185 in185 0 DC -0.800000
v186 in186 0 DC -0.800000
v187 in187 0 DC -0.800000
v188 in188 0 DC -0.800000
v189 in189 0 DC -0.800000
v190 in190 0 DC -0.800000
v191 in191 0 DC -0.800000
v192 in192 0 DC -0.800000
v193 in193 0 DC -0.800000
v194 in194 0 DC -0.800000
v195 in195 0 DC -0.800000
v196 in196 0 DC -0.800000
v197 in197 0 DC -0.800000
v198 in198 0 DC -0.800000
v199 in199 0 DC -0.800000
v200 in200 0 DC -0.800000
v201 in201 0 DC -0.800000
v202 in202 0 DC -0.800000
v203 in203 0 DC -0.800000
v204 in204 0 DC -0.800000
v205 in205 0 DC -0.800000
v206 in206 0 DC -0.109803
v207 in207 0 DC 0.392157
v208 in208 0 DC 0.774902
v209 in209 0 DC 0.774902
v210 in210 0 DC 0.774902
v211 in211 0 DC 0.787451
v212 in212 0 DC 0.260392
v213 in213 0 DC -0.116078
v214 in214 0 DC -0.410981
v215 in215 0 DC -0.800000
v216 in216 0 DC -0.800000
v217 in217 0 DC -0.800000
v218 in218 0 DC -0.800000
v219 in219 0 DC -0.800000
v220 in220 0 DC -0.800000
v221 in221 0 DC -0.800000
v222 in222 0 DC -0.800000
v223 in223 0 DC -0.800000
v224 in224 0 DC -0.800000
v225 in225 0 DC -0.800000
v226 in226 0 DC -0.800000
v227 in227 0 DC -0.800000
v228 in228 0 DC -0.800000
v229 in229 0 DC -0.800000
v230 in230 0 DC -0.800000
v231 in231 0 DC -0.800000
v232 in232 0 DC -0.800000
v233 in233 0 DC -0.800000
v234 in234 0 DC 0.787451
v235 in235 0 DC 0.774902
v236 in236 0 DC 0.774902
v237 in237 0 DC 0.774902
v238 in238 0 DC 0.774902
v239 in239 0 DC 0.787451
v240 in240 0 DC 0.774902
v241 in241 0 DC 0.774902
v242 in242 0 DC 0.580392
v243 in243 0 DC -0.480000
v244 in244 0 DC -0.800000
v245 in245 0 DC -0.800000
v246 in246 0 DC -0.800000
v247 in247 0 DC -0.800000
v248 in248 0 DC -0.800000
v249 in249 0 DC -0.800000
v250 in250 0 DC -0.800000
v251 in251 0 DC -0.800000
v252 in252 0 DC -0.800000
v253 in253 0 DC -0.800000
v254 in254 0 DC -0.800000
v255 in255 0 DC -0.800000
v256 in256 0 DC -0.800000
v257 in257 0 DC -0.800000
v258 in258 0 DC -0.800000
v259 in259 0 DC -0.800000
v260 in260 0 DC -0.800000
v261 in261 0 DC 0.341962
v262 in262 0 DC 0.800000
v263 in263 0 DC 0.787451
v264 in264 0 DC 0.787451
v265 in265 0 DC 0.787451
v266 in266 0 DC 0.787451
v267 in267 0 DC 0.668235
v268 in268 0 DC 0.592941
v269 in269 0 DC 0.787451
v270 in270 0 DC 0.787451
v271 in271 0 DC 0.787451
v272 in272 0 DC -0.800000
v273 in273 0 DC -0.800000
v274 in274 0 DC -0.800000
v275 in275 0 DC -0.800000
v276 in276 0 DC -0.800000
v277 in277 0 DC -0.800000
v278 in278 0 DC -0.800000
v279 in279 0 DC -0.800000
v280 in280 0 DC -0.800000
v281 in281 0 DC -0.800000
v282 in282 0 DC -0.800000
v283 in283 0 DC -0.800000
v284 in284 0 DC -0.800000
v285 in285 0 DC -0.800000
v286 in286 0 DC -0.800000
v287 in287 0 DC -0.800000
v288 in288 0 DC -0.404706
v289 in289 0 DC 0.586667
v290 in290 0 DC 0.787451
v291 in291 0 DC 0.774902
v292 in292 0 DC 0.774902
v293 in293 0 DC 0.774902
v294 in294 0 DC 0.122354
v295 in295 0 DC -0.316862
v296 in296 0 DC -0.410981
v297 in297 0 DC 0.003138
v298 in298 0 DC 0.774902
v299 in299 0 DC 0.774902
v300 in300 0 DC -0.141176
v301 in301 0 DC -0.800000
v302 in302 0 DC -0.800000
v303 in303 0 DC -0.800000
v304 in304 0 DC -0.800000
v305 in305 0 DC -0.800000
v306 in306 0 DC -0.800000
v307 in307 0 DC -0.800000
v308 in308 0 DC -0.800000
v309 in309 0 DC -0.800000
v310 in310 0 DC -0.800000
v311 in311 0 DC -0.800000
v312 in312 0 DC -0.800000
v313 in313 0 DC -0.800000
v314 in314 0 DC -0.800000
v315 in315 0 DC -0.599216
v316 in316 0 DC 0.649411
v317 in317 0 DC 0.774902
v318 in318 0 DC 0.787451
v319 in319 0 DC 0.774902
v320 in320 0 DC 0.580392
v321 in321 0 DC 0.059608
v322 in322 0 DC -0.737254
v323 in323 0 DC -0.800000
v324 in324 0 DC -0.800000
v325 in325 0 DC -0.605490
v326 in326 0 DC 0.643138
v327 in327 0 DC 0.774902
v328 in328 0 DC 0.724706
v329 in329 0 DC -0.090981
v330 in330 0 DC -0.768627
v331 in331 0 DC -0.800000
v332 in332 0 DC -0.800000
v333 in333 0 DC -0.800000
v334 in334 0 DC -0.800000
v335 in335 0 DC -0.800000
v336 in336 0 DC -0.800000
v337 in337 0 DC -0.800000
v338 in338 0 DC -0.800000
v339 in339 0 DC -0.800000
v340 in340 0 DC -0.800000
v341 in341 0 DC -0.800000
v342 in342 0 DC -0.800000
v343 in343 0 DC -0.567843
v344 in344 0 DC 0.774902
v345 in345 0 DC 0.774902
v346 in346 0 DC 0.787451
v347 in347 0 DC 0.379608
v348 in348 0 DC -0.674510
v349 in349 0 DC -0.800000
v350 in350 0 DC -0.800000
v351 in351 0 DC -0.800000
v352 in352 0 DC -0.800000
v353 in353 0 DC -0.800000
v354 in354 0 DC -0.116078
v355 in355 0 DC 0.774902
v356 in356 0 DC 0.787451
v357 in357 0 DC 0.774902
v358 in358 0 DC -0.580392
v359 in359 0 DC -0.800000
v360 in360 0 DC -0.800000
v361 in361 0 DC -0.800000
v362 in362 0 DC -0.800000
v363 in363 0 DC -0.800000
v364 in364 0 DC -0.800000
v365 in365 0 DC -0.800000
v366 in366 0 DC -0.800000
v367 in367 0 DC -0.800000
v368 in368 0 DC -0.800000
v369 in369 0 DC -0.800000
v370 in370 0 DC -0.800000
v371 in371 0 DC -0.567843
v372 in372 0 DC 0.774902
v373 in373 0 DC 0.774902
v374 in374 0 DC 0.461176
v375 in375 0 DC -0.611765
v376 in376 0 DC -0.800000
v377 in377 0 DC -0.800000
v378 in378 0 DC -0.800000
v379 in379 0 DC -0.800000
v380 in380 0 DC -0.800000
v381 in381 0 DC -0.800000
v382 in382 0 DC -0.605490
v383 in383 0 DC 0.454902
v384 in384 0 DC 0.787451
v385 in385 0 DC 0.774902
v386 in386 0 DC -0.580392
v387 in387 0 DC -0.800000
v388 in388 0 DC -0.800000
v389 in389 0 DC -0.800000
v390 in390 0 DC -0.800000
v391 in391 0 DC -0.800000
v392 in392 0 DC -0.800000
v393 in393 0 DC -0.800000
v394 in394 0 DC -0.800000
v395 in395 0 DC -0.800000
v396 in396 0 DC -0.800000
v397 in397 0 DC -0.800000
v398 in398 0 DC -0.800000
v399 in399 0 DC -0.567843
v400 in400 0 DC 0.787451
v401 in401 0 DC 0.787451
v402 in402 0 DC -0.800000
v403 in403 0 DC -0.800000
v404 in404 0 DC -0.800000
v405 in405 0 DC -0.800000
v406 in406 0 DC -0.800000
v407 in407 0 DC -0.800000
v408 in408 0 DC -0.800000
v409 in409 0 DC -0.800000
v410 in410 0 DC -0.599216
v411 in411 0 DC 0.467451
v412 in412 0 DC 0.800000
v413 in413 0 DC 0.787451
v414 in414 0 DC 0.229019
v415 in415 0 DC -0.800000
v416 in416 0 DC -0.800000
v417 in417 0 DC -0.800000
v418 in418 0 DC -0.800000
v419 in419 0 DC -0.800000
v420 in420 0 DC -0.800000
v421 in421 0 DC -0.800000
v422 in422 0 DC -0.800000
v423 in423 0 DC -0.800000
v424 in424 0 DC -0.800000
v425 in425 0 DC -0.800000
v426 in426 0 DC -0.800000
v427 in427 0 DC 0.078432
v428 in428 0 DC 0.774902
v429 in429 0 DC 0.774902
v430 in430 0 DC -0.800000
v431 in431 0 DC -0.800000
v432 in432 0 DC -0.800000
v433 in433 0 DC -0.800000
v434 in434 0 DC -0.800000
v435 in435 0 DC -0.800000
v436 in436 0 DC -0.800000
v437 in437 0 DC -0.800000
v438 in438 0 DC -0.116078
v439 in439 0 DC 0.774902
v440 in440 0 DC 0.787451
v441 in441 0 DC 0.774902
v442 in442 0 DC -0.580392
v443 in443 0 DC -0.800000
v444 in444 0 DC -0.800000
v445 in445 0 DC -0.800000
v446 in446 0 DC -0.800000
v447 in447 0 DC -0.800000
v448 in448 0 DC -0.800000
v449 in449 0 DC -0.800000
v450 in450 0 DC -0.800000
v451 in451 0 DC -0.800000
v452 in452 0 DC -0.800000
v453 in453 0 DC -0.800000
v454 in454 0 DC -0.800000
v455 in455 0 DC 0.561568
v456 in456 0 DC 0.774902
v457 in457 0 DC 0.774902
v458 in458 0 DC -0.800000
v459 in459 0 DC -0.800000
v460 in460 0 DC -0.800000
v461 in461 0 DC -0.800000
v462 in462 0 DC -0.800000
v463 in463 0 DC -0.800000
v464 in464 0 DC -0.668235
v465 in465 0 DC -0.404706
v466 in466 0 DC 0.649411
v467 in467 0 DC 0.774902
v468 in468 0 DC 0.787451
v469 in469 0 DC 0.643138
v470 in470 0 DC -0.611765
v471 in471 0 DC -0.800000
v472 in472 0 DC -0.800000
v473 in473 0 DC -0.800000
v474 in474 0 DC -0.800000
v475 in475 0 DC -0.800000
v476 in476 0 DC -0.800000
v477 in477 0 DC -0.800000
v478 in478 0 DC -0.800000
v479 in479 0 DC -0.800000
v480 in480 0 DC -0.800000
v481 in481 0 DC -0.800000
v482 in482 0 DC -0.800000
v483 in483 0 DC 0.561568
v484 in484 0 DC 0.774902
v485 in485 0 DC 0.774902
v486 in486 0 DC -0.800000
v487 in487 0 DC -0.800000
v488 in488 0 DC -0.800000
v489 in489 0 DC -0.800000
v490 in490 0 DC -0.800000
v491 in491 0 DC -0.800000
v492 in492 0 DC 0.103530
v493 in493 0 DC 0.774902
v494 in494 0 DC 0.774902
v495 in495 0 DC 0.774902
v496 in496 0 DC 0.586667
v497 in497 0 DC -0.417254
v498 in498 0 DC -0.800000
v499 in499 0 DC -0.800000
v500 in500 0 DC -0.800000
v501 in501 0 DC -0.800000
v502 in502 0 DC -0.800000
v503 in503 0 DC -0.800000
v504 in504 0 DC -0.800000
v505 in505 0 DC -0.800000
v506 in506 0 DC -0.800000
v507 in507 0 DC -0.800000
v508 in508 0 DC -0.800000
v509 in509 0 DC -0.800000
v510 in510 0 DC -0.800000
v511 in511 0 DC 0.561568
v512 in512 0 DC 0.774902
v513 in513 0 DC 0.774902
v514 in514 0 DC -0.800000
v515 in515 0 DC -0.800000
v516 in516 0 DC -0.800000
v517 in517 0 DC -0.800000
v518 in518 0 DC -0.800000
v519 in519 0 DC 0.341962
v520 in520 0 DC 0.586667
v521 in521 0 DC 0.774902
v522 in522 0 DC 0.774902
v523 in523 0 DC 0.774902
v524 in524 0 DC 0.329411
v525 in525 0 DC -0.800000
v526 in526 0 DC -0.800000
v527 in527 0 DC -0.800000
v528 in528 0 DC -0.800000
v529 in529 0 DC -0.800000
v530 in530 0 DC -0.800000
v531 in531 0 DC -0.800000
v532 in532 0 DC -0.800000
v533 in533 0 DC -0.800000
v534 in534 0 DC -0.800000
v535 in535 0 DC -0.800000
v536 in536 0 DC -0.800000
v537 in537 0 DC -0.800000
v538 in538 0 DC -0.800000
v539 in539 0 DC 0.567843
v540 in540 0 DC 0.787451
v541 in541 0 DC 0.787451
v542 in542 0 DC -0.341960
v543 in543 0 DC -0.341960
v544 in544 0 DC 0.630589
v545 in545 0 DC 0.787451
v546 in546 0 DC 0.787451
v547 in547 0 DC 0.800000
v548 in548 0 DC 0.787451
v549 in549 0 DC 0.787451
v550 in550 0 DC 0.787451
v551 in551 0 DC 0.787451
v552 in552 0 DC -0.800000
v553 in553 0 DC -0.800000
v554 in554 0 DC -0.800000
v555 in555 0 DC -0.800000
v556 in556 0 DC -0.800000
v557 in557 0 DC -0.800000
v558 in558 0 DC -0.800000
v559 in559 0 DC -0.800000
v560 in560 0 DC -0.800000
v561 in561 0 DC -0.800000
v562 in562 0 DC -0.800000
v563 in563 0 DC -0.800000
v564 in564 0 DC -0.800000
v565 in565 0 DC -0.800000
v566 in566 0 DC -0.800000
v567 in567 0 DC -0.090981
v568 in568 0 DC 0.774902
v569 in569 0 DC 0.774902
v570 in570 0 DC 0.787451
v571 in571 0 DC 0.774902
v572 in572 0 DC 0.774902
v573 in573 0 DC 0.774902
v574 in574 0 DC 0.774902
v575 in575 0 DC 0.787451
v576 in576 0 DC 0.774902
v577 in577 0 DC 0.774902
v578 in578 0 DC 0.774902
v579 in579 0 DC 0.122354
v580 in580 0 DC -0.800000
v581 in581 0 DC -0.800000
v582 in582 0 DC -0.800000
v583 in583 0 DC -0.800000
v584 in584 0 DC -0.800000
v585 in585 0 DC -0.800000
v586 in586 0 DC -0.800000
v587 in587 0 DC -0.800000
v588 in588 0 DC -0.800000
v589 in589 0 DC -0.800000
v590 in590 0 DC -0.800000
v591 in591 0 DC -0.800000
v592 in592 0 DC -0.800000
v593 in593 0 DC -0.800000
v594 in594 0 DC -0.800000
v595 in595 0 DC -0.605490
v596 in596 0 DC 0.643138
v597 in597 0 DC 0.774902
v598 in598 0 DC 0.787451
v599 in599 0 DC 0.774902
v600 in600 0 DC 0.774902
v601 in601 0 DC 0.774902
v602 in602 0 DC 0.774902
v603 in603 0 DC 0.787451
v604 in604 0 DC 0.643138
v605 in605 0 DC 0.385882
v606 in606 0 DC -0.580392
v607 in607 0 DC -0.737254
v608 in608 0 DC -0.800000
v609 in609 0 DC -0.800000
v610 in610 0 DC -0.800000
v611 in611 0 DC -0.800000
v612 in612 0 DC -0.800000
v613 in613 0 DC -0.800000
v614 in614 0 DC -0.800000
v615 in615 0 DC -0.800000
v616 in616 0 DC -0.800000
v617 in617 0 DC -0.800000
v618 in618 0 DC -0.800000
v619 in619 0 DC -0.800000
v620 in620 0 DC -0.800000
v621 in621 0 DC -0.800000
v622 in622 0 DC -0.800000
v623 in623 0 DC -0.800000
v624 in624 0 DC -0.410981
v625 in625 0 DC 0.090981
v626 in626 0 DC 0.787451
v627 in627 0 DC 0.774902
v628 in628 0 DC 0.774902
v629 in629 0 DC 0.774902
v630 in630 0 DC 0.774902
v631 in631 0 DC 0.787451
v632 in632 0 DC -0.128627
v633 in633 0 DC -0.800000
v634 in634 0 DC -0.800000
v635 in635 0 DC -0.800000
v636 in636 0 DC -0.800000
v637 in637 0 DC -0.800000
v638 in638 0 DC -0.800000
v639 in639 0 DC -0.800000
v640 in640 0 DC -0.800000
v641 in641 0 DC -0.800000
v642 in642 0 DC -0.800000
v643 in643 0 DC -0.800000
v644 in644 0 DC -0.800000
v645 in645 0 DC -0.800000
v646 in646 0 DC -0.800000
v647 in647 0 DC -0.800000
v648 in648 0 DC -0.800000
v649 in649 0 DC -0.800000
v650 in650 0 DC -0.800000
v651 in651 0 DC -0.800000
v652 in652 0 DC -0.800000
v653 in653 0 DC -0.800000
v654 in654 0 DC -0.348235
v655 in655 0 DC 0.291765
v656 in656 0 DC 0.774902
v657 in657 0 DC 0.285490
v658 in658 0 DC -0.354510
v659 in659 0 DC -0.348235
v660 in660 0 DC -0.611765
v661 in661 0 DC -0.800000
v662 in662 0 DC -0.800000
v663 in663 0 DC -0.800000
v664 in664 0 DC -0.800000
v665 in665 0 DC -0.800000
v666 in666 0 DC -0.800000
v667 in667 0 DC -0.800000
v668 in668 0 DC -0.800000
v669 in669 0 DC -0.800000
v670 in670 0 DC -0.800000
v671 in671 0 DC -0.800000
v672 in672 0 DC -0.800000
v673 in673 0 DC -0.800000
v674 in674 0 DC -0.800000
v675 in675 0 DC -0.800000
v676 in676 0 DC -0.800000
v677 in677 0 DC -0.800000
v678 in678 0 DC -0.800000
v679 in679 0 DC -0.800000
v680 in680 0 DC -0.800000
v681 in681 0 DC -0.800000
v682 in682 0 DC -0.800000
v683 in683 0 DC -0.800000
v684 in684 0 DC -0.800000
v685 in685 0 DC -0.800000
v686 in686 0 DC -0.800000
v687 in687 0 DC -0.800000
v688 in688 0 DC -0.800000
v689 in689 0 DC -0.800000
v690 in690 0 DC -0.800000
v691 in691 0 DC -0.800000
v692 in692 0 DC -0.800000
v693 in693 0 DC -0.800000
v694 in694 0 DC -0.800000
v695 in695 0 DC -0.800000
v696 in696 0 DC -0.800000
v697 in697 0 DC -0.800000
v698 in698 0 DC -0.800000
v699 in699 0 DC -0.800000
v700 in700 0 DC -0.800000
v701 in701 0 DC -0.800000
v702 in702 0 DC -0.800000
v703 in703 0 DC -0.800000
v704 in704 0 DC -0.800000
v705 in705 0 DC -0.800000
v706 in706 0 DC -0.800000
v707 in707 0 DC -0.800000
v708 in708 0 DC -0.800000
v709 in709 0 DC -0.800000
v710 in710 0 DC -0.800000
v711 in711 0 DC -0.800000
v712 in712 0 DC -0.800000
v713 in713 0 DC -0.800000
v714 in714 0 DC -0.800000
v715 in715 0 DC -0.800000
v716 in716 0 DC -0.800000
v717 in717 0 DC -0.800000
v718 in718 0 DC -0.800000
v719 in719 0 DC -0.800000
v720 in720 0 DC -0.800000
v721 in721 0 DC -0.800000
v722 in722 0 DC -0.800000
v723 in723 0 DC -0.800000
v724 in724 0 DC -0.800000
v725 in725 0 DC -0.800000
v726 in726 0 DC -0.800000
v727 in727 0 DC -0.800000
v728 in728 0 DC -0.800000
v729 in729 0 DC -0.800000
v730 in730 0 DC -0.800000
v731 in731 0 DC -0.800000
v732 in732 0 DC -0.800000
v733 in733 0 DC -0.800000
v734 in734 0 DC -0.800000
v735 in735 0 DC -0.800000
v736 in736 0 DC -0.800000
v737 in737 0 DC -0.800000
v738 in738 0 DC -0.800000
v739 in739 0 DC -0.800000
v740 in740 0 DC -0.800000
v741 in741 0 DC -0.800000
v742 in742 0 DC -0.800000
v743 in743 0 DC -0.800000
v744 in744 0 DC -0.800000
v745 in745 0 DC -0.800000
v746 in746 0 DC -0.800000
v747 in747 0 DC -0.800000
v748 in748 0 DC -0.800000
v749 in749 0 DC -0.800000
v750 in750 0 DC -0.800000
v751 in751 0 DC -0.800000
v752 in752 0 DC -0.800000
v753 in753 0 DC -0.800000
v754 in754 0 DC -0.800000
v755 in755 0 DC -0.800000
v756 in756 0 DC -0.800000
v757 in757 0 DC -0.800000
v758 in758 0 DC -0.800000
v759 in759 0 DC -0.800000
v760 in760 0 DC -0.800000
v761 in761 0 DC -0.800000
v762 in762 0 DC -0.800000
v763 in763 0 DC -0.800000
v764 in764 0 DC -0.800000
v765 in765 0 DC -0.800000
v766 in766 0 DC -0.800000
v767 in767 0 DC -0.800000
v768 in768 0 DC -0.800000
v769 in769 0 DC -0.800000
v770 in770 0 DC -0.800000
v771 in771 0 DC -0.800000
v772 in772 0 DC -0.800000
v773 in773 0 DC -0.800000
v774 in774 0 DC -0.800000
v775 in775 0 DC -0.800000
v776 in776 0 DC -0.800000
v777 in777 0 DC -0.800000
v778 in778 0 DC -0.800000
v779 in779 0 DC -0.800000
v780 in780 0 DC -0.800000
v781 in781 0 DC -0.800000
v782 in782 0 DC -0.800000
v783 in783 0 DC -0.800000



vss vss 0 DC VssVal



vdd vdd 0 DC VddVal
.TRAN 0.1n tsampling
.MEASURE TRAN pwr AVG 'i(vdd)*VddVal' FROM=0n TO=tsampling
.MEASURE TRAN powr AVG POWER FROM=0n TO=tsampling
.MEAS TRAN VOUT0 FIND v(output0) AT=tsampling
.MEAS TRAN VOUT1 FIND v(output1) AT=tsampling
.MEAS TRAN VOUT2 FIND v(output2) AT=tsampling
.MEAS TRAN VOUT3 FIND v(output3) AT=tsampling
.MEAS TRAN VOUT4 FIND v(output4) AT=tsampling
.MEAS TRAN VOUT5 FIND v(output5) AT=tsampling
.MEAS TRAN VOUT6 FIND v(output6) AT=tsampling
.MEAS TRAN VOUT7 FIND v(output7) AT=tsampling
.MEAS TRAN VOUT8 FIND v(output8) AT=tsampling
.MEAS TRAN VOUT9 FIND v(output9) AT=tsampling

.SUBCKT layer2 vdd vss in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15 in16 in17 in18 in19 in20 in21 in22 in23 in24 in25 in26 in27 in28 in29 in30 in31 in32 in33 in34 in35 in36 in37 in38 in39 in40 in41 in42 in43 in44 in45 in46 in47 in48 in49 in50 in51 in52 in53 in54 in55 in56 in57 in58 in59 in60 in61 in62 in63 in64 in65 in66 in67 in68 in69 in70 in71 in72 in73 in74 in75 in76 in77 in78 in79 in80 in81 in82 in83 in84 in85 in86 in87 in88 in89 in90 in91 in92 in93 in94 in95 in96 in97 in98 in99 in100 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 

**********Non-Negative Weighted Array****************
Rwpos1_1 in1 sp1 22281692032865348.000000
Rwpos1_2 in1 sp2 22281692032865348.000000
Rwpos1_3 in1 sp3 22281692032865348.000000
Rwpos1_4 in1 sp4 21220659078919380.000000
Rwpos1_5 in1 sp5 21220659078919380.000000
Rwpos1_6 in1 sp6 21220659078919380.000000
Rwpos1_7 in1 sp7 21220659078919380.000000
Rwpos1_8 in1 sp8 22281692032865348.000000
Rwpos1_9 in1 sp9 21220659078919380.000000
Rwpos1_10 in1 sp10 21220659078919380.000000
Rwpos2_1 in2 sp1 21220659078919380.000000
Rwpos2_2 in2 sp2 21220659078919380.000000
Rwpos2_3 in2 sp3 21220659078919380.000000
Rwpos2_4 in2 sp4 21220659078919380.000000
Rwpos2_5 in2 sp5 21220659078919380.000000
Rwpos2_6 in2 sp6 22281692032865348.000000
Rwpos2_7 in2 sp7 21220659078919380.000000
Rwpos2_8 in2 sp8 21220659078919380.000000
Rwpos2_9 in2 sp9 22281692032865348.000000
Rwpos2_10 in2 sp10 21220659078919380.000000
Rwpos3_1 in3 sp1 21220659078919380.000000
Rwpos3_2 in3 sp2 21220659078919380.000000
Rwpos3_3 in3 sp3 21220659078919380.000000
Rwpos3_4 in3 sp4 22281692032865348.000000
Rwpos3_5 in3 sp5 21220659078919380.000000
Rwpos3_6 in3 sp6 22281692032865348.000000
Rwpos3_7 in3 sp7 21220659078919380.000000
Rwpos3_8 in3 sp8 22281692032865348.000000
Rwpos3_9 in3 sp9 21220659078919380.000000
Rwpos3_10 in3 sp10 21220659078919380.000000
Rwpos4_1 in4 sp1 22281692032865348.000000
Rwpos4_2 in4 sp2 21220659078919380.000000
Rwpos4_3 in4 sp3 21220659078919380.000000
Rwpos4_4 in4 sp4 21220659078919380.000000
Rwpos4_5 in4 sp5 21220659078919380.000000
Rwpos4_6 in4 sp6 22281692032865348.000000
Rwpos4_7 in4 sp7 21220659078919380.000000
Rwpos4_8 in4 sp8 22281692032865348.000000
Rwpos4_9 in4 sp9 22281692032865348.000000
Rwpos4_10 in4 sp10 21220659078919380.000000
Rwpos5_1 in5 sp1 22281692032865348.000000
Rwpos5_2 in5 sp2 21220659078919380.000000
Rwpos5_3 in5 sp3 21220659078919380.000000
Rwpos5_4 in5 sp4 21220659078919380.000000
Rwpos5_5 in5 sp5 21220659078919380.000000
Rwpos5_6 in5 sp6 22281692032865348.000000
Rwpos5_7 in5 sp7 22281692032865348.000000
Rwpos5_8 in5 sp8 21220659078919380.000000
Rwpos5_9 in5 sp9 21220659078919380.000000
Rwpos5_10 in5 sp10 21220659078919380.000000
Rwpos6_1 in6 sp1 21220659078919380.000000
Rwpos6_2 in6 sp2 22281692032865348.000000
Rwpos6_3 in6 sp3 21220659078919380.000000
Rwpos6_4 in6 sp4 22281692032865348.000000
Rwpos6_5 in6 sp5 22281692032865348.000000
Rwpos6_6 in6 sp6 21220659078919380.000000
Rwpos6_7 in6 sp7 21220659078919380.000000
Rwpos6_8 in6 sp8 21220659078919380.000000
Rwpos6_9 in6 sp9 21220659078919380.000000
Rwpos6_10 in6 sp10 21220659078919380.000000
Rwpos7_1 in7 sp1 21220659078919380.000000
Rwpos7_2 in7 sp2 21220659078919380.000000
Rwpos7_3 in7 sp3 22281692032865348.000000
Rwpos7_4 in7 sp4 22281692032865348.000000
Rwpos7_5 in7 sp5 21220659078919380.000000
Rwpos7_6 in7 sp6 21220659078919380.000000
Rwpos7_7 in7 sp7 21220659078919380.000000
Rwpos7_8 in7 sp8 21220659078919380.000000
Rwpos7_9 in7 sp9 21220659078919380.000000
Rwpos7_10 in7 sp10 22281692032865348.000000
Rwpos8_1 in8 sp1 21220659078919380.000000
Rwpos8_2 in8 sp2 22281692032865348.000000
Rwpos8_3 in8 sp3 22281692032865348.000000
Rwpos8_4 in8 sp4 21220659078919380.000000
Rwpos8_5 in8 sp5 21220659078919380.000000
Rwpos8_6 in8 sp6 21220659078919380.000000
Rwpos8_7 in8 sp7 22281692032865348.000000
Rwpos8_8 in8 sp8 22281692032865348.000000
Rwpos8_9 in8 sp9 22281692032865348.000000
Rwpos8_10 in8 sp10 21220659078919380.000000
Rwpos9_1 in9 sp1 22281692032865348.000000
Rwpos9_2 in9 sp2 21220659078919380.000000
Rwpos9_3 in9 sp3 21220659078919380.000000
Rwpos9_4 in9 sp4 21220659078919380.000000
Rwpos9_5 in9 sp5 22281692032865348.000000
Rwpos9_6 in9 sp6 21220659078919380.000000
Rwpos9_7 in9 sp7 22281692032865348.000000
Rwpos9_8 in9 sp8 21220659078919380.000000
Rwpos9_9 in9 sp9 22281692032865348.000000
Rwpos9_10 in9 sp10 21220659078919380.000000
Rwpos10_1 in10 sp1 21220659078919380.000000
Rwpos10_2 in10 sp2 21220659078919380.000000
Rwpos10_3 in10 sp3 21220659078919380.000000
Rwpos10_4 in10 sp4 21220659078919380.000000
Rwpos10_5 in10 sp5 22281692032865348.000000
Rwpos10_6 in10 sp6 22281692032865348.000000
Rwpos10_7 in10 sp7 21220659078919380.000000
Rwpos10_8 in10 sp8 22281692032865348.000000
Rwpos10_9 in10 sp9 21220659078919380.000000
Rwpos10_10 in10 sp10 21220659078919380.000000
Rwpos11_1 in11 sp1 22281692032865348.000000
Rwpos11_2 in11 sp2 21220659078919380.000000
Rwpos11_3 in11 sp3 21220659078919380.000000
Rwpos11_4 in11 sp4 21220659078919380.000000
Rwpos11_5 in11 sp5 21220659078919380.000000
Rwpos11_6 in11 sp6 21220659078919380.000000
Rwpos11_7 in11 sp7 21220659078919380.000000
Rwpos11_8 in11 sp8 22281692032865348.000000
Rwpos11_9 in11 sp9 21220659078919380.000000
Rwpos11_10 in11 sp10 22281692032865348.000000
Rwpos12_1 in12 sp1 21220659078919380.000000
Rwpos12_2 in12 sp2 21220659078919380.000000
Rwpos12_3 in12 sp3 21220659078919380.000000
Rwpos12_4 in12 sp4 22281692032865348.000000
Rwpos12_5 in12 sp5 21220659078919380.000000
Rwpos12_6 in12 sp6 22281692032865348.000000
Rwpos12_7 in12 sp7 21220659078919380.000000
Rwpos12_8 in12 sp8 22281692032865348.000000
Rwpos12_9 in12 sp9 21220659078919380.000000
Rwpos12_10 in12 sp10 21220659078919380.000000
Rwpos13_1 in13 sp1 21220659078919380.000000
Rwpos13_2 in13 sp2 21220659078919380.000000
Rwpos13_3 in13 sp3 21220659078919380.000000
Rwpos13_4 in13 sp4 21220659078919380.000000
Rwpos13_5 in13 sp5 21220659078919380.000000
Rwpos13_6 in13 sp6 22281692032865348.000000
Rwpos13_7 in13 sp7 21220659078919380.000000
Rwpos13_8 in13 sp8 21220659078919380.000000
Rwpos13_9 in13 sp9 21220659078919380.000000
Rwpos13_10 in13 sp10 22281692032865348.000000
Rwpos14_1 in14 sp1 22281692032865348.000000
Rwpos14_2 in14 sp2 22281692032865348.000000
Rwpos14_3 in14 sp3 21220659078919380.000000
Rwpos14_4 in14 sp4 21220659078919380.000000
Rwpos14_5 in14 sp5 22281692032865348.000000
Rwpos14_6 in14 sp6 21220659078919380.000000
Rwpos14_7 in14 sp7 22281692032865348.000000
Rwpos14_8 in14 sp8 22281692032865348.000000
Rwpos14_9 in14 sp9 21220659078919380.000000
Rwpos14_10 in14 sp10 21220659078919380.000000
Rwpos15_1 in15 sp1 21220659078919380.000000
Rwpos15_2 in15 sp2 22281692032865348.000000
Rwpos15_3 in15 sp3 21220659078919380.000000
Rwpos15_4 in15 sp4 21220659078919380.000000
Rwpos15_5 in15 sp5 21220659078919380.000000
Rwpos15_6 in15 sp6 21220659078919380.000000
Rwpos15_7 in15 sp7 21220659078919380.000000
Rwpos15_8 in15 sp8 21220659078919380.000000
Rwpos15_9 in15 sp9 21220659078919380.000000
Rwpos15_10 in15 sp10 22281692032865348.000000
Rwpos16_1 in16 sp1 22281692032865348.000000
Rwpos16_2 in16 sp2 22281692032865348.000000
Rwpos16_3 in16 sp3 22281692032865348.000000
Rwpos16_4 in16 sp4 22281692032865348.000000
Rwpos16_5 in16 sp5 21220659078919380.000000
Rwpos16_6 in16 sp6 21220659078919380.000000
Rwpos16_7 in16 sp7 21220659078919380.000000
Rwpos16_8 in16 sp8 21220659078919380.000000
Rwpos16_9 in16 sp9 21220659078919380.000000
Rwpos16_10 in16 sp10 22281692032865348.000000
Rwpos17_1 in17 sp1 21220659078919380.000000
Rwpos17_2 in17 sp2 22281692032865348.000000
Rwpos17_3 in17 sp3 21220659078919380.000000
Rwpos17_4 in17 sp4 22281692032865348.000000
Rwpos17_5 in17 sp5 22281692032865348.000000
Rwpos17_6 in17 sp6 21220659078919380.000000
Rwpos17_7 in17 sp7 21220659078919380.000000
Rwpos17_8 in17 sp8 21220659078919380.000000
Rwpos17_9 in17 sp9 22281692032865348.000000
Rwpos17_10 in17 sp10 21220659078919380.000000
Rwpos18_1 in18 sp1 22281692032865348.000000
Rwpos18_2 in18 sp2 21220659078919380.000000
Rwpos18_3 in18 sp3 21220659078919380.000000
Rwpos18_4 in18 sp4 21220659078919380.000000
Rwpos18_5 in18 sp5 21220659078919380.000000
Rwpos18_6 in18 sp6 22281692032865348.000000
Rwpos18_7 in18 sp7 22281692032865348.000000
Rwpos18_8 in18 sp8 21220659078919380.000000
Rwpos18_9 in18 sp9 21220659078919380.000000
Rwpos18_10 in18 sp10 22281692032865348.000000
Rwpos19_1 in19 sp1 21220659078919380.000000
Rwpos19_2 in19 sp2 21220659078919380.000000
Rwpos19_3 in19 sp3 21220659078919380.000000
Rwpos19_4 in19 sp4 22281692032865348.000000
Rwpos19_5 in19 sp5 21220659078919380.000000
Rwpos19_6 in19 sp6 21220659078919380.000000
Rwpos19_7 in19 sp7 21220659078919380.000000
Rwpos19_8 in19 sp8 21220659078919380.000000
Rwpos19_9 in19 sp9 22281692032865348.000000
Rwpos19_10 in19 sp10 22281692032865348.000000
Rwpos20_1 in20 sp1 21220659078919380.000000
Rwpos20_2 in20 sp2 22281692032865348.000000
Rwpos20_3 in20 sp3 21220659078919380.000000
Rwpos20_4 in20 sp4 21220659078919380.000000
Rwpos20_5 in20 sp5 22281692032865348.000000
Rwpos20_6 in20 sp6 22281692032865348.000000
Rwpos20_7 in20 sp7 21220659078919380.000000
Rwpos20_8 in20 sp8 21220659078919380.000000
Rwpos20_9 in20 sp9 22281692032865348.000000
Rwpos20_10 in20 sp10 21220659078919380.000000
Rwpos21_1 in21 sp1 21220659078919380.000000
Rwpos21_2 in21 sp2 21220659078919380.000000
Rwpos21_3 in21 sp3 22281692032865348.000000
Rwpos21_4 in21 sp4 21220659078919380.000000
Rwpos21_5 in21 sp5 22281692032865348.000000
Rwpos21_6 in21 sp6 22281692032865348.000000
Rwpos21_7 in21 sp7 21220659078919380.000000
Rwpos21_8 in21 sp8 22281692032865348.000000
Rwpos21_9 in21 sp9 21220659078919380.000000
Rwpos21_10 in21 sp10 21220659078919380.000000
Rwpos22_1 in22 sp1 21220659078919380.000000
Rwpos22_2 in22 sp2 22281692032865348.000000
Rwpos22_3 in22 sp3 21220659078919380.000000
Rwpos22_4 in22 sp4 22281692032865348.000000
Rwpos22_5 in22 sp5 22281692032865348.000000
Rwpos22_6 in22 sp6 21220659078919380.000000
Rwpos22_7 in22 sp7 21220659078919380.000000
Rwpos22_8 in22 sp8 22281692032865348.000000
Rwpos22_9 in22 sp9 21220659078919380.000000
Rwpos22_10 in22 sp10 21220659078919380.000000
Rwpos23_1 in23 sp1 21220659078919380.000000
Rwpos23_2 in23 sp2 22281692032865348.000000
Rwpos23_3 in23 sp3 21220659078919380.000000
Rwpos23_4 in23 sp4 22281692032865348.000000
Rwpos23_5 in23 sp5 21220659078919380.000000
Rwpos23_6 in23 sp6 22281692032865348.000000
Rwpos23_7 in23 sp7 21220659078919380.000000
Rwpos23_8 in23 sp8 22281692032865348.000000
Rwpos23_9 in23 sp9 21220659078919380.000000
Rwpos23_10 in23 sp10 21220659078919380.000000
Rwpos24_1 in24 sp1 21220659078919380.000000
Rwpos24_2 in24 sp2 22281692032865348.000000
Rwpos24_3 in24 sp3 21220659078919380.000000
Rwpos24_4 in24 sp4 21220659078919380.000000
Rwpos24_5 in24 sp5 22281692032865348.000000
Rwpos24_6 in24 sp6 21220659078919380.000000
Rwpos24_7 in24 sp7 22281692032865348.000000
Rwpos24_8 in24 sp8 22281692032865348.000000
Rwpos24_9 in24 sp9 22281692032865348.000000
Rwpos24_10 in24 sp10 21220659078919380.000000
Rwpos25_1 in25 sp1 21220659078919380.000000
Rwpos25_2 in25 sp2 21220659078919380.000000
Rwpos25_3 in25 sp3 22281692032865348.000000
Rwpos25_4 in25 sp4 21220659078919380.000000
Rwpos25_5 in25 sp5 22281692032865348.000000
Rwpos25_6 in25 sp6 21220659078919380.000000
Rwpos25_7 in25 sp7 21220659078919380.000000
Rwpos25_8 in25 sp8 21220659078919380.000000
Rwpos25_9 in25 sp9 22281692032865348.000000
Rwpos25_10 in25 sp10 21220659078919380.000000
Rwpos26_1 in26 sp1 22281692032865348.000000
Rwpos26_2 in26 sp2 21220659078919380.000000
Rwpos26_3 in26 sp3 22281692032865348.000000
Rwpos26_4 in26 sp4 22281692032865348.000000
Rwpos26_5 in26 sp5 21220659078919380.000000
Rwpos26_6 in26 sp6 21220659078919380.000000
Rwpos26_7 in26 sp7 21220659078919380.000000
Rwpos26_8 in26 sp8 22281692032865348.000000
Rwpos26_9 in26 sp9 21220659078919380.000000
Rwpos26_10 in26 sp10 22281692032865348.000000
Rwpos27_1 in27 sp1 21220659078919380.000000
Rwpos27_2 in27 sp2 21220659078919380.000000
Rwpos27_3 in27 sp3 21220659078919380.000000
Rwpos27_4 in27 sp4 21220659078919380.000000
Rwpos27_5 in27 sp5 21220659078919380.000000
Rwpos27_6 in27 sp6 21220659078919380.000000
Rwpos27_7 in27 sp7 22281692032865348.000000
Rwpos27_8 in27 sp8 22281692032865348.000000
Rwpos27_9 in27 sp9 22281692032865348.000000
Rwpos27_10 in27 sp10 22281692032865348.000000
Rwpos28_1 in28 sp1 21220659078919380.000000
Rwpos28_2 in28 sp2 22281692032865348.000000
Rwpos28_3 in28 sp3 21220659078919380.000000
Rwpos28_4 in28 sp4 22281692032865348.000000
Rwpos28_5 in28 sp5 21220659078919380.000000
Rwpos28_6 in28 sp6 22281692032865348.000000
Rwpos28_7 in28 sp7 21220659078919380.000000
Rwpos28_8 in28 sp8 21220659078919380.000000
Rwpos28_9 in28 sp9 21220659078919380.000000
Rwpos28_10 in28 sp10 22281692032865348.000000
Rwpos29_1 in29 sp1 21220659078919380.000000
Rwpos29_2 in29 sp2 21220659078919380.000000
Rwpos29_3 in29 sp3 21220659078919380.000000
Rwpos29_4 in29 sp4 22281692032865348.000000
Rwpos29_5 in29 sp5 21220659078919380.000000
Rwpos29_6 in29 sp6 21220659078919380.000000
Rwpos29_7 in29 sp7 21220659078919380.000000
Rwpos29_8 in29 sp8 22281692032865348.000000
Rwpos29_9 in29 sp9 21220659078919380.000000
Rwpos29_10 in29 sp10 21220659078919380.000000
Rwpos30_1 in30 sp1 22281692032865348.000000
Rwpos30_2 in30 sp2 22281692032865348.000000
Rwpos30_3 in30 sp3 22281692032865348.000000
Rwpos30_4 in30 sp4 21220659078919380.000000
Rwpos30_5 in30 sp5 22281692032865348.000000
Rwpos30_6 in30 sp6 22281692032865348.000000
Rwpos30_7 in30 sp7 21220659078919380.000000
Rwpos30_8 in30 sp8 21220659078919380.000000
Rwpos30_9 in30 sp9 21220659078919380.000000
Rwpos30_10 in30 sp10 21220659078919380.000000
Rwpos31_1 in31 sp1 21220659078919380.000000
Rwpos31_2 in31 sp2 21220659078919380.000000
Rwpos31_3 in31 sp3 22281692032865348.000000
Rwpos31_4 in31 sp4 21220659078919380.000000
Rwpos31_5 in31 sp5 21220659078919380.000000
Rwpos31_6 in31 sp6 21220659078919380.000000
Rwpos31_7 in31 sp7 21220659078919380.000000
Rwpos31_8 in31 sp8 22281692032865348.000000
Rwpos31_9 in31 sp9 22281692032865348.000000
Rwpos31_10 in31 sp10 21220659078919380.000000
Rwpos32_1 in32 sp1 22281692032865348.000000
Rwpos32_2 in32 sp2 21220659078919380.000000
Rwpos32_3 in32 sp3 21220659078919380.000000
Rwpos32_4 in32 sp4 21220659078919380.000000
Rwpos32_5 in32 sp5 22281692032865348.000000
Rwpos32_6 in32 sp6 21220659078919380.000000
Rwpos32_7 in32 sp7 21220659078919380.000000
Rwpos32_8 in32 sp8 21220659078919380.000000
Rwpos32_9 in32 sp9 22281692032865348.000000
Rwpos32_10 in32 sp10 22281692032865348.000000
Rwpos33_1 in33 sp1 21220659078919380.000000
Rwpos33_2 in33 sp2 21220659078919380.000000
Rwpos33_3 in33 sp3 22281692032865348.000000
Rwpos33_4 in33 sp4 22281692032865348.000000
Rwpos33_5 in33 sp5 21220659078919380.000000
Rwpos33_6 in33 sp6 21220659078919380.000000
Rwpos33_7 in33 sp7 21220659078919380.000000
Rwpos33_8 in33 sp8 21220659078919380.000000
Rwpos33_9 in33 sp9 22281692032865348.000000
Rwpos33_10 in33 sp10 21220659078919380.000000
Rwpos34_1 in34 sp1 21220659078919380.000000
Rwpos34_2 in34 sp2 22281692032865348.000000
Rwpos34_3 in34 sp3 21220659078919380.000000
Rwpos34_4 in34 sp4 21220659078919380.000000
Rwpos34_5 in34 sp5 21220659078919380.000000
Rwpos34_6 in34 sp6 21220659078919380.000000
Rwpos34_7 in34 sp7 21220659078919380.000000
Rwpos34_8 in34 sp8 22281692032865348.000000
Rwpos34_9 in34 sp9 21220659078919380.000000
Rwpos34_10 in34 sp10 22281692032865348.000000
Rwpos35_1 in35 sp1 21220659078919380.000000
Rwpos35_2 in35 sp2 22281692032865348.000000
Rwpos35_3 in35 sp3 21220659078919380.000000
Rwpos35_4 in35 sp4 22281692032865348.000000
Rwpos35_5 in35 sp5 21220659078919380.000000
Rwpos35_6 in35 sp6 22281692032865348.000000
Rwpos35_7 in35 sp7 22281692032865348.000000
Rwpos35_8 in35 sp8 21220659078919380.000000
Rwpos35_9 in35 sp9 21220659078919380.000000
Rwpos35_10 in35 sp10 21220659078919380.000000
Rwpos36_1 in36 sp1 21220659078919380.000000
Rwpos36_2 in36 sp2 21220659078919380.000000
Rwpos36_3 in36 sp3 21220659078919380.000000
Rwpos36_4 in36 sp4 22281692032865348.000000
Rwpos36_5 in36 sp5 21220659078919380.000000
Rwpos36_6 in36 sp6 22281692032865348.000000
Rwpos36_7 in36 sp7 22281692032865348.000000
Rwpos36_8 in36 sp8 21220659078919380.000000
Rwpos36_9 in36 sp9 21220659078919380.000000
Rwpos36_10 in36 sp10 21220659078919380.000000
Rwpos37_1 in37 sp1 21220659078919380.000000
Rwpos37_2 in37 sp2 21220659078919380.000000
Rwpos37_3 in37 sp3 21220659078919380.000000
Rwpos37_4 in37 sp4 21220659078919380.000000
Rwpos37_5 in37 sp5 21220659078919380.000000
Rwpos37_6 in37 sp6 21220659078919380.000000
Rwpos37_7 in37 sp7 21220659078919380.000000
Rwpos37_8 in37 sp8 22281692032865348.000000
Rwpos37_9 in37 sp9 21220659078919380.000000
Rwpos37_10 in37 sp10 22281692032865348.000000
Rwpos38_1 in38 sp1 22281692032865348.000000
Rwpos38_2 in38 sp2 22281692032865348.000000
Rwpos38_3 in38 sp3 22281692032865348.000000
Rwpos38_4 in38 sp4 22281692032865348.000000
Rwpos38_5 in38 sp5 21220659078919380.000000
Rwpos38_6 in38 sp6 21220659078919380.000000
Rwpos38_7 in38 sp7 21220659078919380.000000
Rwpos38_8 in38 sp8 21220659078919380.000000
Rwpos38_9 in38 sp9 21220659078919380.000000
Rwpos38_10 in38 sp10 21220659078919380.000000
Rwpos39_1 in39 sp1 21220659078919380.000000
Rwpos39_2 in39 sp2 22281692032865348.000000
Rwpos39_3 in39 sp3 22281692032865348.000000
Rwpos39_4 in39 sp4 21220659078919380.000000
Rwpos39_5 in39 sp5 21220659078919380.000000
Rwpos39_6 in39 sp6 21220659078919380.000000
Rwpos39_7 in39 sp7 21220659078919380.000000
Rwpos39_8 in39 sp8 22281692032865348.000000
Rwpos39_9 in39 sp9 22281692032865348.000000
Rwpos39_10 in39 sp10 21220659078919380.000000
Rwpos40_1 in40 sp1 21220659078919380.000000
Rwpos40_2 in40 sp2 21220659078919380.000000
Rwpos40_3 in40 sp3 22281692032865348.000000
Rwpos40_4 in40 sp4 21220659078919380.000000
Rwpos40_5 in40 sp5 21220659078919380.000000
Rwpos40_6 in40 sp6 21220659078919380.000000
Rwpos40_7 in40 sp7 22281692032865348.000000
Rwpos40_8 in40 sp8 21220659078919380.000000
Rwpos40_9 in40 sp9 21220659078919380.000000
Rwpos40_10 in40 sp10 21220659078919380.000000
Rwpos41_1 in41 sp1 21220659078919380.000000
Rwpos41_2 in41 sp2 21220659078919380.000000
Rwpos41_3 in41 sp3 21220659078919380.000000
Rwpos41_4 in41 sp4 21220659078919380.000000
Rwpos41_5 in41 sp5 21220659078919380.000000
Rwpos41_6 in41 sp6 22281692032865348.000000
Rwpos41_7 in41 sp7 22281692032865348.000000
Rwpos41_8 in41 sp8 21220659078919380.000000
Rwpos41_9 in41 sp9 22281692032865348.000000
Rwpos41_10 in41 sp10 22281692032865348.000000
Rwpos42_1 in42 sp1 21220659078919380.000000
Rwpos42_2 in42 sp2 21220659078919380.000000
Rwpos42_3 in42 sp3 21220659078919380.000000
Rwpos42_4 in42 sp4 22281692032865348.000000
Rwpos42_5 in42 sp5 22281692032865348.000000
Rwpos42_6 in42 sp6 21220659078919380.000000
Rwpos42_7 in42 sp7 22281692032865348.000000
Rwpos42_8 in42 sp8 21220659078919380.000000
Rwpos42_9 in42 sp9 21220659078919380.000000
Rwpos42_10 in42 sp10 21220659078919380.000000
Rwpos43_1 in43 sp1 21220659078919380.000000
Rwpos43_2 in43 sp2 21220659078919380.000000
Rwpos43_3 in43 sp3 21220659078919380.000000
Rwpos43_4 in43 sp4 22281692032865348.000000
Rwpos43_5 in43 sp5 22281692032865348.000000
Rwpos43_6 in43 sp6 21220659078919380.000000
Rwpos43_7 in43 sp7 22281692032865348.000000
Rwpos43_8 in43 sp8 22281692032865348.000000
Rwpos43_9 in43 sp9 21220659078919380.000000
Rwpos43_10 in43 sp10 21220659078919380.000000
Rwpos44_1 in44 sp1 22281692032865348.000000
Rwpos44_2 in44 sp2 21220659078919380.000000
Rwpos44_3 in44 sp3 21220659078919380.000000
Rwpos44_4 in44 sp4 21220659078919380.000000
Rwpos44_5 in44 sp5 21220659078919380.000000
Rwpos44_6 in44 sp6 21220659078919380.000000
Rwpos44_7 in44 sp7 22281692032865348.000000
Rwpos44_8 in44 sp8 22281692032865348.000000
Rwpos44_9 in44 sp9 21220659078919380.000000
Rwpos44_10 in44 sp10 22281692032865348.000000
Rwpos45_1 in45 sp1 21220659078919380.000000
Rwpos45_2 in45 sp2 21220659078919380.000000
Rwpos45_3 in45 sp3 22281692032865348.000000
Rwpos45_4 in45 sp4 22281692032865348.000000
Rwpos45_5 in45 sp5 21220659078919380.000000
Rwpos45_6 in45 sp6 22281692032865348.000000
Rwpos45_7 in45 sp7 21220659078919380.000000
Rwpos45_8 in45 sp8 21220659078919380.000000
Rwpos45_9 in45 sp9 21220659078919380.000000
Rwpos45_10 in45 sp10 21220659078919380.000000
Rwpos46_1 in46 sp1 21220659078919380.000000
Rwpos46_2 in46 sp2 21220659078919380.000000
Rwpos46_3 in46 sp3 22281692032865348.000000
Rwpos46_4 in46 sp4 21220659078919380.000000
Rwpos46_5 in46 sp5 21220659078919380.000000
Rwpos46_6 in46 sp6 22281692032865348.000000
Rwpos46_7 in46 sp7 22281692032865348.000000
Rwpos46_8 in46 sp8 21220659078919380.000000
Rwpos46_9 in46 sp9 21220659078919380.000000
Rwpos46_10 in46 sp10 22281692032865348.000000
Rwpos47_1 in47 sp1 22281692032865348.000000
Rwpos47_2 in47 sp2 21220659078919380.000000
Rwpos47_3 in47 sp3 22281692032865348.000000
Rwpos47_4 in47 sp4 22281692032865348.000000
Rwpos47_5 in47 sp5 21220659078919380.000000
Rwpos47_6 in47 sp6 21220659078919380.000000
Rwpos47_7 in47 sp7 21220659078919380.000000
Rwpos47_8 in47 sp8 22281692032865348.000000
Rwpos47_9 in47 sp9 22281692032865348.000000
Rwpos47_10 in47 sp10 21220659078919380.000000
Rwpos48_1 in48 sp1 21220659078919380.000000
Rwpos48_2 in48 sp2 22281692032865348.000000
Rwpos48_3 in48 sp3 21220659078919380.000000
Rwpos48_4 in48 sp4 21220659078919380.000000
Rwpos48_5 in48 sp5 22281692032865348.000000
Rwpos48_6 in48 sp6 21220659078919380.000000
Rwpos48_7 in48 sp7 22281692032865348.000000
Rwpos48_8 in48 sp8 21220659078919380.000000
Rwpos48_9 in48 sp9 21220659078919380.000000
Rwpos48_10 in48 sp10 21220659078919380.000000
Rwpos49_1 in49 sp1 22281692032865348.000000
Rwpos49_2 in49 sp2 21220659078919380.000000
Rwpos49_3 in49 sp3 21220659078919380.000000
Rwpos49_4 in49 sp4 21220659078919380.000000
Rwpos49_5 in49 sp5 21220659078919380.000000
Rwpos49_6 in49 sp6 22281692032865348.000000
Rwpos49_7 in49 sp7 22281692032865348.000000
Rwpos49_8 in49 sp8 21220659078919380.000000
Rwpos49_9 in49 sp9 21220659078919380.000000
Rwpos49_10 in49 sp10 21220659078919380.000000
Rwpos50_1 in50 sp1 21220659078919380.000000
Rwpos50_2 in50 sp2 22281692032865348.000000
Rwpos50_3 in50 sp3 21220659078919380.000000
Rwpos50_4 in50 sp4 21220659078919380.000000
Rwpos50_5 in50 sp5 21220659078919380.000000
Rwpos50_6 in50 sp6 21220659078919380.000000
Rwpos50_7 in50 sp7 22281692032865348.000000
Rwpos50_8 in50 sp8 21220659078919380.000000
Rwpos50_9 in50 sp9 21220659078919380.000000
Rwpos50_10 in50 sp10 22281692032865348.000000
Rwpos51_1 in51 sp1 22281692032865348.000000
Rwpos51_2 in51 sp2 21220659078919380.000000
Rwpos51_3 in51 sp3 21220659078919380.000000
Rwpos51_4 in51 sp4 22281692032865348.000000
Rwpos51_5 in51 sp5 21220659078919380.000000
Rwpos51_6 in51 sp6 21220659078919380.000000
Rwpos51_7 in51 sp7 21220659078919380.000000
Rwpos51_8 in51 sp8 22281692032865348.000000
Rwpos51_9 in51 sp9 21220659078919380.000000
Rwpos51_10 in51 sp10 21220659078919380.000000
Rwpos52_1 in52 sp1 21220659078919380.000000
Rwpos52_2 in52 sp2 21220659078919380.000000
Rwpos52_3 in52 sp3 22281692032865348.000000
Rwpos52_4 in52 sp4 21220659078919380.000000
Rwpos52_5 in52 sp5 21220659078919380.000000
Rwpos52_6 in52 sp6 22281692032865348.000000
Rwpos52_7 in52 sp7 21220659078919380.000000
Rwpos52_8 in52 sp8 22281692032865348.000000
Rwpos52_9 in52 sp9 21220659078919380.000000
Rwpos52_10 in52 sp10 21220659078919380.000000
Rwpos53_1 in53 sp1 21220659078919380.000000
Rwpos53_2 in53 sp2 22281692032865348.000000
Rwpos53_3 in53 sp3 21220659078919380.000000
Rwpos53_4 in53 sp4 21220659078919380.000000
Rwpos53_5 in53 sp5 22281692032865348.000000
Rwpos53_6 in53 sp6 21220659078919380.000000
Rwpos53_7 in53 sp7 21220659078919380.000000
Rwpos53_8 in53 sp8 22281692032865348.000000
Rwpos53_9 in53 sp9 21220659078919380.000000
Rwpos53_10 in53 sp10 22281692032865348.000000
Rwpos54_1 in54 sp1 21220659078919380.000000
Rwpos54_2 in54 sp2 21220659078919380.000000
Rwpos54_3 in54 sp3 22281692032865348.000000
Rwpos54_4 in54 sp4 22281692032865348.000000
Rwpos54_5 in54 sp5 21220659078919380.000000
Rwpos54_6 in54 sp6 22281692032865348.000000
Rwpos54_7 in54 sp7 21220659078919380.000000
Rwpos54_8 in54 sp8 22281692032865348.000000
Rwpos54_9 in54 sp9 21220659078919380.000000
Rwpos54_10 in54 sp10 21220659078919380.000000
Rwpos55_1 in55 sp1 21220659078919380.000000
Rwpos55_2 in55 sp2 21220659078919380.000000
Rwpos55_3 in55 sp3 21220659078919380.000000
Rwpos55_4 in55 sp4 21220659078919380.000000
Rwpos55_5 in55 sp5 21220659078919380.000000
Rwpos55_6 in55 sp6 22281692032865348.000000
Rwpos55_7 in55 sp7 21220659078919380.000000
Rwpos55_8 in55 sp8 21220659078919380.000000
Rwpos55_9 in55 sp9 22281692032865348.000000
Rwpos55_10 in55 sp10 22281692032865348.000000
Rwpos56_1 in56 sp1 21220659078919380.000000
Rwpos56_2 in56 sp2 21220659078919380.000000
Rwpos56_3 in56 sp3 22281692032865348.000000
Rwpos56_4 in56 sp4 22281692032865348.000000
Rwpos56_5 in56 sp5 22281692032865348.000000
Rwpos56_6 in56 sp6 22281692032865348.000000
Rwpos56_7 in56 sp7 21220659078919380.000000
Rwpos56_8 in56 sp8 22281692032865348.000000
Rwpos56_9 in56 sp9 21220659078919380.000000
Rwpos56_10 in56 sp10 21220659078919380.000000
Rwpos57_1 in57 sp1 21220659078919380.000000
Rwpos57_2 in57 sp2 21220659078919380.000000
Rwpos57_3 in57 sp3 22281692032865348.000000
Rwpos57_4 in57 sp4 21220659078919380.000000
Rwpos57_5 in57 sp5 21220659078919380.000000
Rwpos57_6 in57 sp6 21220659078919380.000000
Rwpos57_7 in57 sp7 21220659078919380.000000
Rwpos57_8 in57 sp8 21220659078919380.000000
Rwpos57_9 in57 sp9 22281692032865348.000000
Rwpos57_10 in57 sp10 22281692032865348.000000
Rwpos58_1 in58 sp1 21220659078919380.000000
Rwpos58_2 in58 sp2 21220659078919380.000000
Rwpos58_3 in58 sp3 22281692032865348.000000
Rwpos58_4 in58 sp4 21220659078919380.000000
Rwpos58_5 in58 sp5 22281692032865348.000000
Rwpos58_6 in58 sp6 21220659078919380.000000
Rwpos58_7 in58 sp7 21220659078919380.000000
Rwpos58_8 in58 sp8 21220659078919380.000000
Rwpos58_9 in58 sp9 21220659078919380.000000
Rwpos58_10 in58 sp10 22281692032865348.000000
Rwpos59_1 in59 sp1 21220659078919380.000000
Rwpos59_2 in59 sp2 22281692032865348.000000
Rwpos59_3 in59 sp3 22281692032865348.000000
Rwpos59_4 in59 sp4 21220659078919380.000000
Rwpos59_5 in59 sp5 21220659078919380.000000
Rwpos59_6 in59 sp6 22281692032865348.000000
Rwpos59_7 in59 sp7 21220659078919380.000000
Rwpos59_8 in59 sp8 21220659078919380.000000
Rwpos59_9 in59 sp9 21220659078919380.000000
Rwpos59_10 in59 sp10 21220659078919380.000000
Rwpos60_1 in60 sp1 22281692032865348.000000
Rwpos60_2 in60 sp2 22281692032865348.000000
Rwpos60_3 in60 sp3 21220659078919380.000000
Rwpos60_4 in60 sp4 21220659078919380.000000
Rwpos60_5 in60 sp5 21220659078919380.000000
Rwpos60_6 in60 sp6 21220659078919380.000000
Rwpos60_7 in60 sp7 22281692032865348.000000
Rwpos60_8 in60 sp8 21220659078919380.000000
Rwpos60_9 in60 sp9 21220659078919380.000000
Rwpos60_10 in60 sp10 21220659078919380.000000
Rwpos61_1 in61 sp1 21220659078919380.000000
Rwpos61_2 in61 sp2 21220659078919380.000000
Rwpos61_3 in61 sp3 21220659078919380.000000
Rwpos61_4 in61 sp4 21220659078919380.000000
Rwpos61_5 in61 sp5 22281692032865348.000000
Rwpos61_6 in61 sp6 22281692032865348.000000
Rwpos61_7 in61 sp7 21220659078919380.000000
Rwpos61_8 in61 sp8 22281692032865348.000000
Rwpos61_9 in61 sp9 22281692032865348.000000
Rwpos61_10 in61 sp10 21220659078919380.000000
Rwpos62_1 in62 sp1 21220659078919380.000000
Rwpos62_2 in62 sp2 22281692032865348.000000
Rwpos62_3 in62 sp3 22281692032865348.000000
Rwpos62_4 in62 sp4 21220659078919380.000000
Rwpos62_5 in62 sp5 21220659078919380.000000
Rwpos62_6 in62 sp6 21220659078919380.000000
Rwpos62_7 in62 sp7 22281692032865348.000000
Rwpos62_8 in62 sp8 22281692032865348.000000
Rwpos62_9 in62 sp9 22281692032865348.000000
Rwpos62_10 in62 sp10 21220659078919380.000000
Rwpos63_1 in63 sp1 21220659078919380.000000
Rwpos63_2 in63 sp2 22281692032865348.000000
Rwpos63_3 in63 sp3 21220659078919380.000000
Rwpos63_4 in63 sp4 21220659078919380.000000
Rwpos63_5 in63 sp5 21220659078919380.000000
Rwpos63_6 in63 sp6 22281692032865348.000000
Rwpos63_7 in63 sp7 22281692032865348.000000
Rwpos63_8 in63 sp8 22281692032865348.000000
Rwpos63_9 in63 sp9 21220659078919380.000000
Rwpos63_10 in63 sp10 21220659078919380.000000
Rwpos64_1 in64 sp1 21220659078919380.000000
Rwpos64_2 in64 sp2 21220659078919380.000000
Rwpos64_3 in64 sp3 21220659078919380.000000
Rwpos64_4 in64 sp4 21220659078919380.000000
Rwpos64_5 in64 sp5 22281692032865348.000000
Rwpos64_6 in64 sp6 21220659078919380.000000
Rwpos64_7 in64 sp7 21220659078919380.000000
Rwpos64_8 in64 sp8 21220659078919380.000000
Rwpos64_9 in64 sp9 21220659078919380.000000
Rwpos64_10 in64 sp10 21220659078919380.000000
Rwpos65_1 in65 sp1 22281692032865348.000000
Rwpos65_2 in65 sp2 21220659078919380.000000
Rwpos65_3 in65 sp3 22281692032865348.000000
Rwpos65_4 in65 sp4 21220659078919380.000000
Rwpos65_5 in65 sp5 21220659078919380.000000
Rwpos65_6 in65 sp6 21220659078919380.000000
Rwpos65_7 in65 sp7 21220659078919380.000000
Rwpos65_8 in65 sp8 21220659078919380.000000
Rwpos65_9 in65 sp9 22281692032865348.000000
Rwpos65_10 in65 sp10 21220659078919380.000000
Rwpos66_1 in66 sp1 21220659078919380.000000
Rwpos66_2 in66 sp2 22281692032865348.000000
Rwpos66_3 in66 sp3 21220659078919380.000000
Rwpos66_4 in66 sp4 22281692032865348.000000
Rwpos66_5 in66 sp5 22281692032865348.000000
Rwpos66_6 in66 sp6 21220659078919380.000000
Rwpos66_7 in66 sp7 21220659078919380.000000
Rwpos66_8 in66 sp8 22281692032865348.000000
Rwpos66_9 in66 sp9 21220659078919380.000000
Rwpos66_10 in66 sp10 21220659078919380.000000
Rwpos67_1 in67 sp1 21220659078919380.000000
Rwpos67_2 in67 sp2 21220659078919380.000000
Rwpos67_3 in67 sp3 22281692032865348.000000
Rwpos67_4 in67 sp4 21220659078919380.000000
Rwpos67_5 in67 sp5 21220659078919380.000000
Rwpos67_6 in67 sp6 22281692032865348.000000
Rwpos67_7 in67 sp7 22281692032865348.000000
Rwpos67_8 in67 sp8 21220659078919380.000000
Rwpos67_9 in67 sp9 21220659078919380.000000
Rwpos67_10 in67 sp10 21220659078919380.000000
Rwpos68_1 in68 sp1 22281692032865348.000000
Rwpos68_2 in68 sp2 21220659078919380.000000
Rwpos68_3 in68 sp3 21220659078919380.000000
Rwpos68_4 in68 sp4 21220659078919380.000000
Rwpos68_5 in68 sp5 21220659078919380.000000
Rwpos68_6 in68 sp6 22281692032865348.000000
Rwpos68_7 in68 sp7 21220659078919380.000000
Rwpos68_8 in68 sp8 21220659078919380.000000
Rwpos68_9 in68 sp9 21220659078919380.000000
Rwpos68_10 in68 sp10 21220659078919380.000000
Rwpos69_1 in69 sp1 21220659078919380.000000
Rwpos69_2 in69 sp2 22281692032865348.000000
Rwpos69_3 in69 sp3 21220659078919380.000000
Rwpos69_4 in69 sp4 22281692032865348.000000
Rwpos69_5 in69 sp5 21220659078919380.000000
Rwpos69_6 in69 sp6 21220659078919380.000000
Rwpos69_7 in69 sp7 21220659078919380.000000
Rwpos69_8 in69 sp8 21220659078919380.000000
Rwpos69_9 in69 sp9 22281692032865348.000000
Rwpos69_10 in69 sp10 22281692032865348.000000
Rwpos70_1 in70 sp1 21220659078919380.000000
Rwpos70_2 in70 sp2 22281692032865348.000000
Rwpos70_3 in70 sp3 22281692032865348.000000
Rwpos70_4 in70 sp4 21220659078919380.000000
Rwpos70_5 in70 sp5 22281692032865348.000000
Rwpos70_6 in70 sp6 21220659078919380.000000
Rwpos70_7 in70 sp7 21220659078919380.000000
Rwpos70_8 in70 sp8 22281692032865348.000000
Rwpos70_9 in70 sp9 21220659078919380.000000
Rwpos70_10 in70 sp10 21220659078919380.000000
Rwpos71_1 in71 sp1 21220659078919380.000000
Rwpos71_2 in71 sp2 22281692032865348.000000
Rwpos71_3 in71 sp3 22281692032865348.000000
Rwpos71_4 in71 sp4 22281692032865348.000000
Rwpos71_5 in71 sp5 21220659078919380.000000
Rwpos71_6 in71 sp6 22281692032865348.000000
Rwpos71_7 in71 sp7 21220659078919380.000000
Rwpos71_8 in71 sp8 21220659078919380.000000
Rwpos71_9 in71 sp9 21220659078919380.000000
Rwpos71_10 in71 sp10 22281692032865348.000000
Rwpos72_1 in72 sp1 21220659078919380.000000
Rwpos72_2 in72 sp2 21220659078919380.000000
Rwpos72_3 in72 sp3 22281692032865348.000000
Rwpos72_4 in72 sp4 22281692032865348.000000
Rwpos72_5 in72 sp5 22281692032865348.000000
Rwpos72_6 in72 sp6 21220659078919380.000000
Rwpos72_7 in72 sp7 21220659078919380.000000
Rwpos72_8 in72 sp8 21220659078919380.000000
Rwpos72_9 in72 sp9 21220659078919380.000000
Rwpos72_10 in72 sp10 21220659078919380.000000
Rwpos73_1 in73 sp1 22281692032865348.000000
Rwpos73_2 in73 sp2 21220659078919380.000000
Rwpos73_3 in73 sp3 21220659078919380.000000
Rwpos73_4 in73 sp4 22281692032865348.000000
Rwpos73_5 in73 sp5 21220659078919380.000000
Rwpos73_6 in73 sp6 21220659078919380.000000
Rwpos73_7 in73 sp7 21220659078919380.000000
Rwpos73_8 in73 sp8 21220659078919380.000000
Rwpos73_9 in73 sp9 22281692032865348.000000
Rwpos73_10 in73 sp10 22281692032865348.000000
Rwpos74_1 in74 sp1 21220659078919380.000000
Rwpos74_2 in74 sp2 21220659078919380.000000
Rwpos74_3 in74 sp3 21220659078919380.000000
Rwpos74_4 in74 sp4 21220659078919380.000000
Rwpos74_5 in74 sp5 22281692032865348.000000
Rwpos74_6 in74 sp6 22281692032865348.000000
Rwpos74_7 in74 sp7 21220659078919380.000000
Rwpos74_8 in74 sp8 21220659078919380.000000
Rwpos74_9 in74 sp9 21220659078919380.000000
Rwpos74_10 in74 sp10 21220659078919380.000000
Rwpos75_1 in75 sp1 21220659078919380.000000
Rwpos75_2 in75 sp2 21220659078919380.000000
Rwpos75_3 in75 sp3 21220659078919380.000000
Rwpos75_4 in75 sp4 22281692032865348.000000
Rwpos75_5 in75 sp5 21220659078919380.000000
Rwpos75_6 in75 sp6 21220659078919380.000000
Rwpos75_7 in75 sp7 21220659078919380.000000
Rwpos75_8 in75 sp8 22281692032865348.000000
Rwpos75_9 in75 sp9 21220659078919380.000000
Rwpos75_10 in75 sp10 21220659078919380.000000
Rwpos76_1 in76 sp1 21220659078919380.000000
Rwpos76_2 in76 sp2 22281692032865348.000000
Rwpos76_3 in76 sp3 22281692032865348.000000
Rwpos76_4 in76 sp4 22281692032865348.000000
Rwpos76_5 in76 sp5 21220659078919380.000000
Rwpos76_6 in76 sp6 21220659078919380.000000
Rwpos76_7 in76 sp7 21220659078919380.000000
Rwpos76_8 in76 sp8 21220659078919380.000000
Rwpos76_9 in76 sp9 21220659078919380.000000
Rwpos76_10 in76 sp10 22281692032865348.000000
Rwpos77_1 in77 sp1 21220659078919380.000000
Rwpos77_2 in77 sp2 21220659078919380.000000
Rwpos77_3 in77 sp3 22281692032865348.000000
Rwpos77_4 in77 sp4 21220659078919380.000000
Rwpos77_5 in77 sp5 22281692032865348.000000
Rwpos77_6 in77 sp6 21220659078919380.000000
Rwpos77_7 in77 sp7 22281692032865348.000000
Rwpos77_8 in77 sp8 21220659078919380.000000
Rwpos77_9 in77 sp9 21220659078919380.000000
Rwpos77_10 in77 sp10 21220659078919380.000000
Rwpos78_1 in78 sp1 21220659078919380.000000
Rwpos78_2 in78 sp2 21220659078919380.000000
Rwpos78_3 in78 sp3 22281692032865348.000000
Rwpos78_4 in78 sp4 21220659078919380.000000
Rwpos78_5 in78 sp5 21220659078919380.000000
Rwpos78_6 in78 sp6 22281692032865348.000000
Rwpos78_7 in78 sp7 21220659078919380.000000
Rwpos78_8 in78 sp8 21220659078919380.000000
Rwpos78_9 in78 sp9 21220659078919380.000000
Rwpos78_10 in78 sp10 22281692032865348.000000
Rwpos79_1 in79 sp1 21220659078919380.000000
Rwpos79_2 in79 sp2 22281692032865348.000000
Rwpos79_3 in79 sp3 22281692032865348.000000
Rwpos79_4 in79 sp4 21220659078919380.000000
Rwpos79_5 in79 sp5 22281692032865348.000000
Rwpos79_6 in79 sp6 22281692032865348.000000
Rwpos79_7 in79 sp7 21220659078919380.000000
Rwpos79_8 in79 sp8 21220659078919380.000000
Rwpos79_9 in79 sp9 21220659078919380.000000
Rwpos79_10 in79 sp10 21220659078919380.000000
Rwpos80_1 in80 sp1 21220659078919380.000000
Rwpos80_2 in80 sp2 22281692032865348.000000
Rwpos80_3 in80 sp3 21220659078919380.000000
Rwpos80_4 in80 sp4 22281692032865348.000000
Rwpos80_5 in80 sp5 21220659078919380.000000
Rwpos80_6 in80 sp6 22281692032865348.000000
Rwpos80_7 in80 sp7 22281692032865348.000000
Rwpos80_8 in80 sp8 21220659078919380.000000
Rwpos80_9 in80 sp9 21220659078919380.000000
Rwpos80_10 in80 sp10 21220659078919380.000000
Rwpos81_1 in81 sp1 22281692032865348.000000
Rwpos81_2 in81 sp2 22281692032865348.000000
Rwpos81_3 in81 sp3 21220659078919380.000000
Rwpos81_4 in81 sp4 22281692032865348.000000
Rwpos81_5 in81 sp5 21220659078919380.000000
Rwpos81_6 in81 sp6 21220659078919380.000000
Rwpos81_7 in81 sp7 22281692032865348.000000
Rwpos81_8 in81 sp8 22281692032865348.000000
Rwpos81_9 in81 sp9 21220659078919380.000000
Rwpos81_10 in81 sp10 21220659078919380.000000
Rwpos82_1 in82 sp1 22281692032865348.000000
Rwpos82_2 in82 sp2 21220659078919380.000000
Rwpos82_3 in82 sp3 22281692032865348.000000
Rwpos82_4 in82 sp4 21220659078919380.000000
Rwpos82_5 in82 sp5 21220659078919380.000000
Rwpos82_6 in82 sp6 21220659078919380.000000
Rwpos82_7 in82 sp7 22281692032865348.000000
Rwpos82_8 in82 sp8 21220659078919380.000000
Rwpos82_9 in82 sp9 21220659078919380.000000
Rwpos82_10 in82 sp10 21220659078919380.000000
Rwpos83_1 in83 sp1 21220659078919380.000000
Rwpos83_2 in83 sp2 22281692032865348.000000
Rwpos83_3 in83 sp3 22281692032865348.000000
Rwpos83_4 in83 sp4 21220659078919380.000000
Rwpos83_5 in83 sp5 21220659078919380.000000
Rwpos83_6 in83 sp6 21220659078919380.000000
Rwpos83_7 in83 sp7 22281692032865348.000000
Rwpos83_8 in83 sp8 21220659078919380.000000
Rwpos83_9 in83 sp9 21220659078919380.000000
Rwpos83_10 in83 sp10 21220659078919380.000000
Rwpos84_1 in84 sp1 22281692032865348.000000
Rwpos84_2 in84 sp2 21220659078919380.000000
Rwpos84_3 in84 sp3 21220659078919380.000000
Rwpos84_4 in84 sp4 21220659078919380.000000
Rwpos84_5 in84 sp5 22281692032865348.000000
Rwpos84_6 in84 sp6 21220659078919380.000000
Rwpos84_7 in84 sp7 21220659078919380.000000
Rwpos84_8 in84 sp8 21220659078919380.000000
Rwpos84_9 in84 sp9 21220659078919380.000000
Rwpos84_10 in84 sp10 22281692032865348.000000
Rwpos85_1 in85 sp1 22281692032865348.000000
Rwpos85_2 in85 sp2 22281692032865348.000000
Rwpos85_3 in85 sp3 22281692032865348.000000
Rwpos85_4 in85 sp4 21220659078919380.000000
Rwpos85_5 in85 sp5 21220659078919380.000000
Rwpos85_6 in85 sp6 21220659078919380.000000
Rwpos85_7 in85 sp7 22281692032865348.000000
Rwpos85_8 in85 sp8 21220659078919380.000000
Rwpos85_9 in85 sp9 21220659078919380.000000
Rwpos85_10 in85 sp10 22281692032865348.000000
Rwpos86_1 in86 sp1 22281692032865348.000000
Rwpos86_2 in86 sp2 22281692032865348.000000
Rwpos86_3 in86 sp3 21220659078919380.000000
Rwpos86_4 in86 sp4 21220659078919380.000000
Rwpos86_5 in86 sp5 22281692032865348.000000
Rwpos86_6 in86 sp6 21220659078919380.000000
Rwpos86_7 in86 sp7 21220659078919380.000000
Rwpos86_8 in86 sp8 21220659078919380.000000
Rwpos86_9 in86 sp9 21220659078919380.000000
Rwpos86_10 in86 sp10 21220659078919380.000000
Rwpos87_1 in87 sp1 21220659078919380.000000
Rwpos87_2 in87 sp2 22281692032865348.000000
Rwpos87_3 in87 sp3 21220659078919380.000000
Rwpos87_4 in87 sp4 21220659078919380.000000
Rwpos87_5 in87 sp5 21220659078919380.000000
Rwpos87_6 in87 sp6 22281692032865348.000000
Rwpos87_7 in87 sp7 21220659078919380.000000
Rwpos87_8 in87 sp8 21220659078919380.000000
Rwpos87_9 in87 sp9 21220659078919380.000000
Rwpos87_10 in87 sp10 22281692032865348.000000
Rwpos88_1 in88 sp1 21220659078919380.000000
Rwpos88_2 in88 sp2 21220659078919380.000000
Rwpos88_3 in88 sp3 21220659078919380.000000
Rwpos88_4 in88 sp4 21220659078919380.000000
Rwpos88_5 in88 sp5 22281692032865348.000000
Rwpos88_6 in88 sp6 22281692032865348.000000
Rwpos88_7 in88 sp7 21220659078919380.000000
Rwpos88_8 in88 sp8 21220659078919380.000000
Rwpos88_9 in88 sp9 21220659078919380.000000
Rwpos88_10 in88 sp10 22281692032865348.000000
Rwpos89_1 in89 sp1 21220659078919380.000000
Rwpos89_2 in89 sp2 21220659078919380.000000
Rwpos89_3 in89 sp3 22281692032865348.000000
Rwpos89_4 in89 sp4 22281692032865348.000000
Rwpos89_5 in89 sp5 21220659078919380.000000
Rwpos89_6 in89 sp6 21220659078919380.000000
Rwpos89_7 in89 sp7 21220659078919380.000000
Rwpos89_8 in89 sp8 21220659078919380.000000
Rwpos89_9 in89 sp9 21220659078919380.000000
Rwpos89_10 in89 sp10 22281692032865348.000000
Rwpos90_1 in90 sp1 21220659078919380.000000
Rwpos90_2 in90 sp2 21220659078919380.000000
Rwpos90_3 in90 sp3 21220659078919380.000000
Rwpos90_4 in90 sp4 22281692032865348.000000
Rwpos90_5 in90 sp5 21220659078919380.000000
Rwpos90_6 in90 sp6 22281692032865348.000000
Rwpos90_7 in90 sp7 21220659078919380.000000
Rwpos90_8 in90 sp8 21220659078919380.000000
Rwpos90_9 in90 sp9 21220659078919380.000000
Rwpos90_10 in90 sp10 22281692032865348.000000
Rwpos91_1 in91 sp1 21220659078919380.000000
Rwpos91_2 in91 sp2 21220659078919380.000000
Rwpos91_3 in91 sp3 22281692032865348.000000
Rwpos91_4 in91 sp4 21220659078919380.000000
Rwpos91_5 in91 sp5 21220659078919380.000000
Rwpos91_6 in91 sp6 21220659078919380.000000
Rwpos91_7 in91 sp7 22281692032865348.000000
Rwpos91_8 in91 sp8 22281692032865348.000000
Rwpos91_9 in91 sp9 21220659078919380.000000
Rwpos91_10 in91 sp10 21220659078919380.000000
Rwpos92_1 in92 sp1 21220659078919380.000000
Rwpos92_2 in92 sp2 21220659078919380.000000
Rwpos92_3 in92 sp3 21220659078919380.000000
Rwpos92_4 in92 sp4 21220659078919380.000000
Rwpos92_5 in92 sp5 21220659078919380.000000
Rwpos92_6 in92 sp6 21220659078919380.000000
Rwpos92_7 in92 sp7 21220659078919380.000000
Rwpos92_8 in92 sp8 21220659078919380.000000
Rwpos92_9 in92 sp9 21220659078919380.000000
Rwpos92_10 in92 sp10 21220659078919380.000000
Rwpos93_1 in93 sp1 21220659078919380.000000
Rwpos93_2 in93 sp2 22281692032865348.000000
Rwpos93_3 in93 sp3 21220659078919380.000000
Rwpos93_4 in93 sp4 21220659078919380.000000
Rwpos93_5 in93 sp5 21220659078919380.000000
Rwpos93_6 in93 sp6 22281692032865348.000000
Rwpos93_7 in93 sp7 22281692032865348.000000
Rwpos93_8 in93 sp8 22281692032865348.000000
Rwpos93_9 in93 sp9 21220659078919380.000000
Rwpos93_10 in93 sp10 22281692032865348.000000
Rwpos94_1 in94 sp1 21220659078919380.000000
Rwpos94_2 in94 sp2 21220659078919380.000000
Rwpos94_3 in94 sp3 21220659078919380.000000
Rwpos94_4 in94 sp4 21220659078919380.000000
Rwpos94_5 in94 sp5 22281692032865348.000000
Rwpos94_6 in94 sp6 22281692032865348.000000
Rwpos94_7 in94 sp7 21220659078919380.000000
Rwpos94_8 in94 sp8 21220659078919380.000000
Rwpos94_9 in94 sp9 21220659078919380.000000
Rwpos94_10 in94 sp10 22281692032865348.000000
Rwpos95_1 in95 sp1 21220659078919380.000000
Rwpos95_2 in95 sp2 21220659078919380.000000
Rwpos95_3 in95 sp3 21220659078919380.000000
Rwpos95_4 in95 sp4 21220659078919380.000000
Rwpos95_5 in95 sp5 21220659078919380.000000
Rwpos95_6 in95 sp6 22281692032865348.000000
Rwpos95_7 in95 sp7 21220659078919380.000000
Rwpos95_8 in95 sp8 21220659078919380.000000
Rwpos95_9 in95 sp9 22281692032865348.000000
Rwpos95_10 in95 sp10 22281692032865348.000000
Rwpos96_1 in96 sp1 21220659078919380.000000
Rwpos96_2 in96 sp2 21220659078919380.000000
Rwpos96_3 in96 sp3 22281692032865348.000000
Rwpos96_4 in96 sp4 21220659078919380.000000
Rwpos96_5 in96 sp5 22281692032865348.000000
Rwpos96_6 in96 sp6 21220659078919380.000000
Rwpos96_7 in96 sp7 21220659078919380.000000
Rwpos96_8 in96 sp8 21220659078919380.000000
Rwpos96_9 in96 sp9 22281692032865348.000000
Rwpos96_10 in96 sp10 21220659078919380.000000
Rwpos97_1 in97 sp1 21220659078919380.000000
Rwpos97_2 in97 sp2 22281692032865348.000000
Rwpos97_3 in97 sp3 22281692032865348.000000
Rwpos97_4 in97 sp4 21220659078919380.000000
Rwpos97_5 in97 sp5 21220659078919380.000000
Rwpos97_6 in97 sp6 21220659078919380.000000
Rwpos97_7 in97 sp7 21220659078919380.000000
Rwpos97_8 in97 sp8 21220659078919380.000000
Rwpos97_9 in97 sp9 21220659078919380.000000
Rwpos97_10 in97 sp10 21220659078919380.000000
Rwpos98_1 in98 sp1 22281692032865348.000000
Rwpos98_2 in98 sp2 21220659078919380.000000
Rwpos98_3 in98 sp3 21220659078919380.000000
Rwpos98_4 in98 sp4 21220659078919380.000000
Rwpos98_5 in98 sp5 22281692032865348.000000
Rwpos98_6 in98 sp6 21220659078919380.000000
Rwpos98_7 in98 sp7 21220659078919380.000000
Rwpos98_8 in98 sp8 22281692032865348.000000
Rwpos98_9 in98 sp9 21220659078919380.000000
Rwpos98_10 in98 sp10 21220659078919380.000000
Rwpos99_1 in99 sp1 22281692032865348.000000
Rwpos99_2 in99 sp2 22281692032865348.000000
Rwpos99_3 in99 sp3 22281692032865348.000000
Rwpos99_4 in99 sp4 21220659078919380.000000
Rwpos99_5 in99 sp5 22281692032865348.000000
Rwpos99_6 in99 sp6 22281692032865348.000000
Rwpos99_7 in99 sp7 21220659078919380.000000
Rwpos99_8 in99 sp8 21220659078919380.000000
Rwpos99_9 in99 sp9 21220659078919380.000000
Rwpos99_10 in99 sp10 21220659078919380.000000
Rwpos100_1 in100 sp1 21220659078919380.000000
Rwpos100_2 in100 sp2 21220659078919380.000000
Rwpos100_3 in100 sp3 22281692032865348.000000
Rwpos100_4 in100 sp4 21220659078919380.000000
Rwpos100_5 in100 sp5 21220659078919380.000000
Rwpos100_6 in100 sp6 21220659078919380.000000
Rwpos100_7 in100 sp7 21220659078919380.000000
Rwpos100_8 in100 sp8 21220659078919380.000000
Rwpos100_9 in100 sp9 21220659078919380.000000
Rwpos100_10 in100 sp10 21220659078919380.000000


**********Negative Weighted Array****************

Rwneg1_1 in1 sn1 21220659078919380.000000
Rwneg1_2 in1 sn2 21220659078919380.000000
Rwneg1_3 in1 sn3 21220659078919380.000000
Rwneg1_4 in1 sn4 22281692032865348.000000
Rwneg1_5 in1 sn5 22281692032865348.000000
Rwneg1_6 in1 sn6 22281692032865348.000000
Rwneg1_7 in1 sn7 22281692032865348.000000
Rwneg1_8 in1 sn8 21220659078919380.000000
Rwneg1_9 in1 sn9 22281692032865348.000000
Rwneg1_10 in1 sn10 22281692032865348.000000
Rwneg2_1 in2 sn1 21220659078919380.000000
Rwneg2_2 in2 sn2 22281692032865348.000000
Rwneg2_3 in2 sn3 22281692032865348.000000
Rwneg2_4 in2 sn4 21220659078919380.000000
Rwneg2_5 in2 sn5 22281692032865348.000000
Rwneg2_6 in2 sn6 21220659078919380.000000
Rwneg2_7 in2 sn7 22281692032865348.000000
Rwneg2_8 in2 sn8 22281692032865348.000000
Rwneg2_9 in2 sn9 21220659078919380.000000
Rwneg2_10 in2 sn10 22281692032865348.000000
Rwneg3_1 in3 sn1 22281692032865348.000000
Rwneg3_2 in3 sn2 22281692032865348.000000
Rwneg3_3 in3 sn3 22281692032865348.000000
Rwneg3_4 in3 sn4 21220659078919380.000000
Rwneg3_5 in3 sn5 21220659078919380.000000
Rwneg3_6 in3 sn6 21220659078919380.000000
Rwneg3_7 in3 sn7 22281692032865348.000000
Rwneg3_8 in3 sn8 21220659078919380.000000
Rwneg3_9 in3 sn9 22281692032865348.000000
Rwneg3_10 in3 sn10 21220659078919380.000000
Rwneg4_1 in4 sn1 21220659078919380.000000
Rwneg4_2 in4 sn2 22281692032865348.000000
Rwneg4_3 in4 sn3 22281692032865348.000000
Rwneg4_4 in4 sn4 22281692032865348.000000
Rwneg4_5 in4 sn5 22281692032865348.000000
Rwneg4_6 in4 sn6 21220659078919380.000000
Rwneg4_7 in4 sn7 22281692032865348.000000
Rwneg4_8 in4 sn8 21220659078919380.000000
Rwneg4_9 in4 sn9 21220659078919380.000000
Rwneg4_10 in4 sn10 21220659078919380.000000
Rwneg5_1 in5 sn1 21220659078919380.000000
Rwneg5_2 in5 sn2 21220659078919380.000000
Rwneg5_3 in5 sn3 22281692032865348.000000
Rwneg5_4 in5 sn4 22281692032865348.000000
Rwneg5_5 in5 sn5 22281692032865348.000000
Rwneg5_6 in5 sn6 21220659078919380.000000
Rwneg5_7 in5 sn7 21220659078919380.000000
Rwneg5_8 in5 sn8 21220659078919380.000000
Rwneg5_9 in5 sn9 22281692032865348.000000
Rwneg5_10 in5 sn10 22281692032865348.000000
Rwneg6_1 in6 sn1 21220659078919380.000000
Rwneg6_2 in6 sn2 21220659078919380.000000
Rwneg6_3 in6 sn3 21220659078919380.000000
Rwneg6_4 in6 sn4 21220659078919380.000000
Rwneg6_5 in6 sn5 21220659078919380.000000
Rwneg6_6 in6 sn6 22281692032865348.000000
Rwneg6_7 in6 sn7 22281692032865348.000000
Rwneg6_8 in6 sn8 22281692032865348.000000
Rwneg6_9 in6 sn9 22281692032865348.000000
Rwneg6_10 in6 sn10 22281692032865348.000000
Rwneg7_1 in7 sn1 21220659078919380.000000
Rwneg7_2 in7 sn2 21220659078919380.000000
Rwneg7_3 in7 sn3 21220659078919380.000000
Rwneg7_4 in7 sn4 21220659078919380.000000
Rwneg7_5 in7 sn5 22281692032865348.000000
Rwneg7_6 in7 sn6 22281692032865348.000000
Rwneg7_7 in7 sn7 22281692032865348.000000
Rwneg7_8 in7 sn8 22281692032865348.000000
Rwneg7_9 in7 sn9 22281692032865348.000000
Rwneg7_10 in7 sn10 21220659078919380.000000
Rwneg8_1 in8 sn1 22281692032865348.000000
Rwneg8_2 in8 sn2 21220659078919380.000000
Rwneg8_3 in8 sn3 21220659078919380.000000
Rwneg8_4 in8 sn4 22281692032865348.000000
Rwneg8_5 in8 sn5 22281692032865348.000000
Rwneg8_6 in8 sn6 22281692032865348.000000
Rwneg8_7 in8 sn7 21220659078919380.000000
Rwneg8_8 in8 sn8 21220659078919380.000000
Rwneg8_9 in8 sn9 21220659078919380.000000
Rwneg8_10 in8 sn10 22281692032865348.000000
Rwneg9_1 in9 sn1 21220659078919380.000000
Rwneg9_2 in9 sn2 22281692032865348.000000
Rwneg9_3 in9 sn3 22281692032865348.000000
Rwneg9_4 in9 sn4 22281692032865348.000000
Rwneg9_5 in9 sn5 21220659078919380.000000
Rwneg9_6 in9 sn6 22281692032865348.000000
Rwneg9_7 in9 sn7 21220659078919380.000000
Rwneg9_8 in9 sn8 21220659078919380.000000
Rwneg9_9 in9 sn9 21220659078919380.000000
Rwneg9_10 in9 sn10 22281692032865348.000000
Rwneg10_1 in10 sn1 22281692032865348.000000
Rwneg10_2 in10 sn2 22281692032865348.000000
Rwneg10_3 in10 sn3 22281692032865348.000000
Rwneg10_4 in10 sn4 22281692032865348.000000
Rwneg10_5 in10 sn5 21220659078919380.000000
Rwneg10_6 in10 sn6 21220659078919380.000000
Rwneg10_7 in10 sn7 21220659078919380.000000
Rwneg10_8 in10 sn8 21220659078919380.000000
Rwneg10_9 in10 sn9 22281692032865348.000000
Rwneg10_10 in10 sn10 22281692032865348.000000
Rwneg11_1 in11 sn1 21220659078919380.000000
Rwneg11_2 in11 sn2 22281692032865348.000000
Rwneg11_3 in11 sn3 22281692032865348.000000
Rwneg11_4 in11 sn4 22281692032865348.000000
Rwneg11_5 in11 sn5 22281692032865348.000000
Rwneg11_6 in11 sn6 22281692032865348.000000
Rwneg11_7 in11 sn7 22281692032865348.000000
Rwneg11_8 in11 sn8 21220659078919380.000000
Rwneg11_9 in11 sn9 21220659078919380.000000
Rwneg11_10 in11 sn10 21220659078919380.000000
Rwneg12_1 in12 sn1 21220659078919380.000000
Rwneg12_2 in12 sn2 21220659078919380.000000
Rwneg12_3 in12 sn3 22281692032865348.000000
Rwneg12_4 in12 sn4 21220659078919380.000000
Rwneg12_5 in12 sn5 22281692032865348.000000
Rwneg12_6 in12 sn6 21220659078919380.000000
Rwneg12_7 in12 sn7 21220659078919380.000000
Rwneg12_8 in12 sn8 21220659078919380.000000
Rwneg12_9 in12 sn9 22281692032865348.000000
Rwneg12_10 in12 sn10 22281692032865348.000000
Rwneg13_1 in13 sn1 22281692032865348.000000
Rwneg13_2 in13 sn2 22281692032865348.000000
Rwneg13_3 in13 sn3 22281692032865348.000000
Rwneg13_4 in13 sn4 22281692032865348.000000
Rwneg13_5 in13 sn5 22281692032865348.000000
Rwneg13_6 in13 sn6 21220659078919380.000000
Rwneg13_7 in13 sn7 22281692032865348.000000
Rwneg13_8 in13 sn8 22281692032865348.000000
Rwneg13_9 in13 sn9 21220659078919380.000000
Rwneg13_10 in13 sn10 21220659078919380.000000
Rwneg14_1 in14 sn1 21220659078919380.000000
Rwneg14_2 in14 sn2 21220659078919380.000000
Rwneg14_3 in14 sn3 22281692032865348.000000
Rwneg14_4 in14 sn4 22281692032865348.000000
Rwneg14_5 in14 sn5 21220659078919380.000000
Rwneg14_6 in14 sn6 22281692032865348.000000
Rwneg14_7 in14 sn7 21220659078919380.000000
Rwneg14_8 in14 sn8 21220659078919380.000000
Rwneg14_9 in14 sn9 22281692032865348.000000
Rwneg14_10 in14 sn10 22281692032865348.000000
Rwneg15_1 in15 sn1 22281692032865348.000000
Rwneg15_2 in15 sn2 21220659078919380.000000
Rwneg15_3 in15 sn3 22281692032865348.000000
Rwneg15_4 in15 sn4 22281692032865348.000000
Rwneg15_5 in15 sn5 21220659078919380.000000
Rwneg15_6 in15 sn6 22281692032865348.000000
Rwneg15_7 in15 sn7 22281692032865348.000000
Rwneg15_8 in15 sn8 22281692032865348.000000
Rwneg15_9 in15 sn9 22281692032865348.000000
Rwneg15_10 in15 sn10 21220659078919380.000000
Rwneg16_1 in16 sn1 21220659078919380.000000
Rwneg16_2 in16 sn2 21220659078919380.000000
Rwneg16_3 in16 sn3 21220659078919380.000000
Rwneg16_4 in16 sn4 21220659078919380.000000
Rwneg16_5 in16 sn5 22281692032865348.000000
Rwneg16_6 in16 sn6 22281692032865348.000000
Rwneg16_7 in16 sn7 22281692032865348.000000
Rwneg16_8 in16 sn8 22281692032865348.000000
Rwneg16_9 in16 sn9 22281692032865348.000000
Rwneg16_10 in16 sn10 21220659078919380.000000
Rwneg17_1 in17 sn1 22281692032865348.000000
Rwneg17_2 in17 sn2 21220659078919380.000000
Rwneg17_3 in17 sn3 22281692032865348.000000
Rwneg17_4 in17 sn4 21220659078919380.000000
Rwneg17_5 in17 sn5 21220659078919380.000000
Rwneg17_6 in17 sn6 22281692032865348.000000
Rwneg17_7 in17 sn7 22281692032865348.000000
Rwneg17_8 in17 sn8 21220659078919380.000000
Rwneg17_9 in17 sn9 21220659078919380.000000
Rwneg17_10 in17 sn10 22281692032865348.000000
Rwneg18_1 in18 sn1 21220659078919380.000000
Rwneg18_2 in18 sn2 22281692032865348.000000
Rwneg18_3 in18 sn3 22281692032865348.000000
Rwneg18_4 in18 sn4 22281692032865348.000000
Rwneg18_5 in18 sn5 22281692032865348.000000
Rwneg18_6 in18 sn6 21220659078919380.000000
Rwneg18_7 in18 sn7 21220659078919380.000000
Rwneg18_8 in18 sn8 22281692032865348.000000
Rwneg18_9 in18 sn9 21220659078919380.000000
Rwneg18_10 in18 sn10 21220659078919380.000000
Rwneg19_1 in19 sn1 22281692032865348.000000
Rwneg19_2 in19 sn2 22281692032865348.000000
Rwneg19_3 in19 sn3 21220659078919380.000000
Rwneg19_4 in19 sn4 21220659078919380.000000
Rwneg19_5 in19 sn5 22281692032865348.000000
Rwneg19_6 in19 sn6 21220659078919380.000000
Rwneg19_7 in19 sn7 22281692032865348.000000
Rwneg19_8 in19 sn8 22281692032865348.000000
Rwneg19_9 in19 sn9 21220659078919380.000000
Rwneg19_10 in19 sn10 21220659078919380.000000
Rwneg20_1 in20 sn1 22281692032865348.000000
Rwneg20_2 in20 sn2 21220659078919380.000000
Rwneg20_3 in20 sn3 22281692032865348.000000
Rwneg20_4 in20 sn4 22281692032865348.000000
Rwneg20_5 in20 sn5 21220659078919380.000000
Rwneg20_6 in20 sn6 21220659078919380.000000
Rwneg20_7 in20 sn7 22281692032865348.000000
Rwneg20_8 in20 sn8 21220659078919380.000000
Rwneg20_9 in20 sn9 21220659078919380.000000
Rwneg20_10 in20 sn10 22281692032865348.000000
Rwneg21_1 in21 sn1 21220659078919380.000000
Rwneg21_2 in21 sn2 21220659078919380.000000
Rwneg21_3 in21 sn3 21220659078919380.000000
Rwneg21_4 in21 sn4 22281692032865348.000000
Rwneg21_5 in21 sn5 21220659078919380.000000
Rwneg21_6 in21 sn6 21220659078919380.000000
Rwneg21_7 in21 sn7 22281692032865348.000000
Rwneg21_8 in21 sn8 21220659078919380.000000
Rwneg21_9 in21 sn9 22281692032865348.000000
Rwneg21_10 in21 sn10 22281692032865348.000000
Rwneg22_1 in22 sn1 22281692032865348.000000
Rwneg22_2 in22 sn2 21220659078919380.000000
Rwneg22_3 in22 sn3 22281692032865348.000000
Rwneg22_4 in22 sn4 21220659078919380.000000
Rwneg22_5 in22 sn5 21220659078919380.000000
Rwneg22_6 in22 sn6 22281692032865348.000000
Rwneg22_7 in22 sn7 22281692032865348.000000
Rwneg22_8 in22 sn8 21220659078919380.000000
Rwneg22_9 in22 sn9 22281692032865348.000000
Rwneg22_10 in22 sn10 22281692032865348.000000
Rwneg23_1 in23 sn1 22281692032865348.000000
Rwneg23_2 in23 sn2 21220659078919380.000000
Rwneg23_3 in23 sn3 22281692032865348.000000
Rwneg23_4 in23 sn4 21220659078919380.000000
Rwneg23_5 in23 sn5 21220659078919380.000000
Rwneg23_6 in23 sn6 21220659078919380.000000
Rwneg23_7 in23 sn7 21220659078919380.000000
Rwneg23_8 in23 sn8 21220659078919380.000000
Rwneg23_9 in23 sn9 22281692032865348.000000
Rwneg23_10 in23 sn10 22281692032865348.000000
Rwneg24_1 in24 sn1 22281692032865348.000000
Rwneg24_2 in24 sn2 21220659078919380.000000
Rwneg24_3 in24 sn3 22281692032865348.000000
Rwneg24_4 in24 sn4 22281692032865348.000000
Rwneg24_5 in24 sn5 21220659078919380.000000
Rwneg24_6 in24 sn6 22281692032865348.000000
Rwneg24_7 in24 sn7 21220659078919380.000000
Rwneg24_8 in24 sn8 21220659078919380.000000
Rwneg24_9 in24 sn9 21220659078919380.000000
Rwneg24_10 in24 sn10 22281692032865348.000000
Rwneg25_1 in25 sn1 22281692032865348.000000
Rwneg25_2 in25 sn2 21220659078919380.000000
Rwneg25_3 in25 sn3 21220659078919380.000000
Rwneg25_4 in25 sn4 22281692032865348.000000
Rwneg25_5 in25 sn5 21220659078919380.000000
Rwneg25_6 in25 sn6 22281692032865348.000000
Rwneg25_7 in25 sn7 21220659078919380.000000
Rwneg25_8 in25 sn8 22281692032865348.000000
Rwneg25_9 in25 sn9 21220659078919380.000000
Rwneg25_10 in25 sn10 22281692032865348.000000
Rwneg26_1 in26 sn1 21220659078919380.000000
Rwneg26_2 in26 sn2 22281692032865348.000000
Rwneg26_3 in26 sn3 21220659078919380.000000
Rwneg26_4 in26 sn4 21220659078919380.000000
Rwneg26_5 in26 sn5 22281692032865348.000000
Rwneg26_6 in26 sn6 22281692032865348.000000
Rwneg26_7 in26 sn7 22281692032865348.000000
Rwneg26_8 in26 sn8 21220659078919380.000000
Rwneg26_9 in26 sn9 22281692032865348.000000
Rwneg26_10 in26 sn10 21220659078919380.000000
Rwneg27_1 in27 sn1 22281692032865348.000000
Rwneg27_2 in27 sn2 22281692032865348.000000
Rwneg27_3 in27 sn3 22281692032865348.000000
Rwneg27_4 in27 sn4 22281692032865348.000000
Rwneg27_5 in27 sn5 21220659078919380.000000
Rwneg27_6 in27 sn6 22281692032865348.000000
Rwneg27_7 in27 sn7 21220659078919380.000000
Rwneg27_8 in27 sn8 21220659078919380.000000
Rwneg27_9 in27 sn9 21220659078919380.000000
Rwneg27_10 in27 sn10 21220659078919380.000000
Rwneg28_1 in28 sn1 22281692032865348.000000
Rwneg28_2 in28 sn2 21220659078919380.000000
Rwneg28_3 in28 sn3 22281692032865348.000000
Rwneg28_4 in28 sn4 21220659078919380.000000
Rwneg28_5 in28 sn5 21220659078919380.000000
Rwneg28_6 in28 sn6 21220659078919380.000000
Rwneg28_7 in28 sn7 22281692032865348.000000
Rwneg28_8 in28 sn8 22281692032865348.000000
Rwneg28_9 in28 sn9 22281692032865348.000000
Rwneg28_10 in28 sn10 21220659078919380.000000
Rwneg29_1 in29 sn1 22281692032865348.000000
Rwneg29_2 in29 sn2 22281692032865348.000000
Rwneg29_3 in29 sn3 22281692032865348.000000
Rwneg29_4 in29 sn4 21220659078919380.000000
Rwneg29_5 in29 sn5 22281692032865348.000000
Rwneg29_6 in29 sn6 21220659078919380.000000
Rwneg29_7 in29 sn7 22281692032865348.000000
Rwneg29_8 in29 sn8 21220659078919380.000000
Rwneg29_9 in29 sn9 21220659078919380.000000
Rwneg29_10 in29 sn10 22281692032865348.000000
Rwneg30_1 in30 sn1 21220659078919380.000000
Rwneg30_2 in30 sn2 21220659078919380.000000
Rwneg30_3 in30 sn3 21220659078919380.000000
Rwneg30_4 in30 sn4 22281692032865348.000000
Rwneg30_5 in30 sn5 21220659078919380.000000
Rwneg30_6 in30 sn6 21220659078919380.000000
Rwneg30_7 in30 sn7 22281692032865348.000000
Rwneg30_8 in30 sn8 21220659078919380.000000
Rwneg30_9 in30 sn9 22281692032865348.000000
Rwneg30_10 in30 sn10 22281692032865348.000000
Rwneg31_1 in31 sn1 21220659078919380.000000
Rwneg31_2 in31 sn2 22281692032865348.000000
Rwneg31_3 in31 sn3 21220659078919380.000000
Rwneg31_4 in31 sn4 22281692032865348.000000
Rwneg31_5 in31 sn5 22281692032865348.000000
Rwneg31_6 in31 sn6 22281692032865348.000000
Rwneg31_7 in31 sn7 22281692032865348.000000
Rwneg31_8 in31 sn8 21220659078919380.000000
Rwneg31_9 in31 sn9 21220659078919380.000000
Rwneg31_10 in31 sn10 22281692032865348.000000
Rwneg32_1 in32 sn1 21220659078919380.000000
Rwneg32_2 in32 sn2 22281692032865348.000000
Rwneg32_3 in32 sn3 22281692032865348.000000
Rwneg32_4 in32 sn4 21220659078919380.000000
Rwneg32_5 in32 sn5 21220659078919380.000000
Rwneg32_6 in32 sn6 22281692032865348.000000
Rwneg32_7 in32 sn7 22281692032865348.000000
Rwneg32_8 in32 sn8 22281692032865348.000000
Rwneg32_9 in32 sn9 21220659078919380.000000
Rwneg32_10 in32 sn10 21220659078919380.000000
Rwneg33_1 in33 sn1 21220659078919380.000000
Rwneg33_2 in33 sn2 22281692032865348.000000
Rwneg33_3 in33 sn3 21220659078919380.000000
Rwneg33_4 in33 sn4 21220659078919380.000000
Rwneg33_5 in33 sn5 21220659078919380.000000
Rwneg33_6 in33 sn6 22281692032865348.000000
Rwneg33_7 in33 sn7 22281692032865348.000000
Rwneg33_8 in33 sn8 22281692032865348.000000
Rwneg33_9 in33 sn9 21220659078919380.000000
Rwneg33_10 in33 sn10 22281692032865348.000000
Rwneg34_1 in34 sn1 22281692032865348.000000
Rwneg34_2 in34 sn2 21220659078919380.000000
Rwneg34_3 in34 sn3 22281692032865348.000000
Rwneg34_4 in34 sn4 22281692032865348.000000
Rwneg34_5 in34 sn5 21220659078919380.000000
Rwneg34_6 in34 sn6 22281692032865348.000000
Rwneg34_7 in34 sn7 21220659078919380.000000
Rwneg34_8 in34 sn8 21220659078919380.000000
Rwneg34_9 in34 sn9 22281692032865348.000000
Rwneg34_10 in34 sn10 21220659078919380.000000
Rwneg35_1 in35 sn1 21220659078919380.000000
Rwneg35_2 in35 sn2 21220659078919380.000000
Rwneg35_3 in35 sn3 22281692032865348.000000
Rwneg35_4 in35 sn4 21220659078919380.000000
Rwneg35_5 in35 sn5 22281692032865348.000000
Rwneg35_6 in35 sn6 21220659078919380.000000
Rwneg35_7 in35 sn7 21220659078919380.000000
Rwneg35_8 in35 sn8 22281692032865348.000000
Rwneg35_9 in35 sn9 22281692032865348.000000
Rwneg35_10 in35 sn10 22281692032865348.000000
Rwneg36_1 in36 sn1 22281692032865348.000000
Rwneg36_2 in36 sn2 22281692032865348.000000
Rwneg36_3 in36 sn3 22281692032865348.000000
Rwneg36_4 in36 sn4 21220659078919380.000000
Rwneg36_5 in36 sn5 22281692032865348.000000
Rwneg36_6 in36 sn6 21220659078919380.000000
Rwneg36_7 in36 sn7 21220659078919380.000000
Rwneg36_8 in36 sn8 22281692032865348.000000
Rwneg36_9 in36 sn9 21220659078919380.000000
Rwneg36_10 in36 sn10 22281692032865348.000000
Rwneg37_1 in37 sn1 22281692032865348.000000
Rwneg37_2 in37 sn2 22281692032865348.000000
Rwneg37_3 in37 sn3 21220659078919380.000000
Rwneg37_4 in37 sn4 21220659078919380.000000
Rwneg37_5 in37 sn5 22281692032865348.000000
Rwneg37_6 in37 sn6 22281692032865348.000000
Rwneg37_7 in37 sn7 22281692032865348.000000
Rwneg37_8 in37 sn8 21220659078919380.000000
Rwneg37_9 in37 sn9 22281692032865348.000000
Rwneg37_10 in37 sn10 21220659078919380.000000
Rwneg38_1 in38 sn1 21220659078919380.000000
Rwneg38_2 in38 sn2 21220659078919380.000000
Rwneg38_3 in38 sn3 21220659078919380.000000
Rwneg38_4 in38 sn4 21220659078919380.000000
Rwneg38_5 in38 sn5 22281692032865348.000000
Rwneg38_6 in38 sn6 22281692032865348.000000
Rwneg38_7 in38 sn7 22281692032865348.000000
Rwneg38_8 in38 sn8 22281692032865348.000000
Rwneg38_9 in38 sn9 22281692032865348.000000
Rwneg38_10 in38 sn10 22281692032865348.000000
Rwneg39_1 in39 sn1 22281692032865348.000000
Rwneg39_2 in39 sn2 21220659078919380.000000
Rwneg39_3 in39 sn3 21220659078919380.000000
Rwneg39_4 in39 sn4 22281692032865348.000000
Rwneg39_5 in39 sn5 22281692032865348.000000
Rwneg39_6 in39 sn6 22281692032865348.000000
Rwneg39_7 in39 sn7 21220659078919380.000000
Rwneg39_8 in39 sn8 21220659078919380.000000
Rwneg39_9 in39 sn9 21220659078919380.000000
Rwneg39_10 in39 sn10 22281692032865348.000000
Rwneg40_1 in40 sn1 22281692032865348.000000
Rwneg40_2 in40 sn2 22281692032865348.000000
Rwneg40_3 in40 sn3 21220659078919380.000000
Rwneg40_4 in40 sn4 21220659078919380.000000
Rwneg40_5 in40 sn5 22281692032865348.000000
Rwneg40_6 in40 sn6 22281692032865348.000000
Rwneg40_7 in40 sn7 21220659078919380.000000
Rwneg40_8 in40 sn8 22281692032865348.000000
Rwneg40_9 in40 sn9 22281692032865348.000000
Rwneg40_10 in40 sn10 22281692032865348.000000
Rwneg41_1 in41 sn1 22281692032865348.000000
Rwneg41_2 in41 sn2 22281692032865348.000000
Rwneg41_3 in41 sn3 22281692032865348.000000
Rwneg41_4 in41 sn4 22281692032865348.000000
Rwneg41_5 in41 sn5 21220659078919380.000000
Rwneg41_6 in41 sn6 21220659078919380.000000
Rwneg41_7 in41 sn7 21220659078919380.000000
Rwneg41_8 in41 sn8 22281692032865348.000000
Rwneg41_9 in41 sn9 21220659078919380.000000
Rwneg41_10 in41 sn10 21220659078919380.000000
Rwneg42_1 in42 sn1 21220659078919380.000000
Rwneg42_2 in42 sn2 22281692032865348.000000
Rwneg42_3 in42 sn3 22281692032865348.000000
Rwneg42_4 in42 sn4 21220659078919380.000000
Rwneg42_5 in42 sn5 21220659078919380.000000
Rwneg42_6 in42 sn6 22281692032865348.000000
Rwneg42_7 in42 sn7 21220659078919380.000000
Rwneg42_8 in42 sn8 22281692032865348.000000
Rwneg42_9 in42 sn9 21220659078919380.000000
Rwneg42_10 in42 sn10 22281692032865348.000000
Rwneg43_1 in43 sn1 22281692032865348.000000
Rwneg43_2 in43 sn2 22281692032865348.000000
Rwneg43_3 in43 sn3 22281692032865348.000000
Rwneg43_4 in43 sn4 21220659078919380.000000
Rwneg43_5 in43 sn5 21220659078919380.000000
Rwneg43_6 in43 sn6 21220659078919380.000000
Rwneg43_7 in43 sn7 21220659078919380.000000
Rwneg43_8 in43 sn8 21220659078919380.000000
Rwneg43_9 in43 sn9 22281692032865348.000000
Rwneg43_10 in43 sn10 22281692032865348.000000
Rwneg44_1 in44 sn1 21220659078919380.000000
Rwneg44_2 in44 sn2 21220659078919380.000000
Rwneg44_3 in44 sn3 22281692032865348.000000
Rwneg44_4 in44 sn4 22281692032865348.000000
Rwneg44_5 in44 sn5 22281692032865348.000000
Rwneg44_6 in44 sn6 21220659078919380.000000
Rwneg44_7 in44 sn7 21220659078919380.000000
Rwneg44_8 in44 sn8 21220659078919380.000000
Rwneg44_9 in44 sn9 22281692032865348.000000
Rwneg44_10 in44 sn10 21220659078919380.000000
Rwneg45_1 in45 sn1 21220659078919380.000000
Rwneg45_2 in45 sn2 22281692032865348.000000
Rwneg45_3 in45 sn3 21220659078919380.000000
Rwneg45_4 in45 sn4 21220659078919380.000000
Rwneg45_5 in45 sn5 22281692032865348.000000
Rwneg45_6 in45 sn6 21220659078919380.000000
Rwneg45_7 in45 sn7 22281692032865348.000000
Rwneg45_8 in45 sn8 22281692032865348.000000
Rwneg45_9 in45 sn9 22281692032865348.000000
Rwneg45_10 in45 sn10 22281692032865348.000000
Rwneg46_1 in46 sn1 22281692032865348.000000
Rwneg46_2 in46 sn2 22281692032865348.000000
Rwneg46_3 in46 sn3 21220659078919380.000000
Rwneg46_4 in46 sn4 22281692032865348.000000
Rwneg46_5 in46 sn5 22281692032865348.000000
Rwneg46_6 in46 sn6 21220659078919380.000000
Rwneg46_7 in46 sn7 21220659078919380.000000
Rwneg46_8 in46 sn8 22281692032865348.000000
Rwneg46_9 in46 sn9 22281692032865348.000000
Rwneg46_10 in46 sn10 21220659078919380.000000
Rwneg47_1 in47 sn1 21220659078919380.000000
Rwneg47_2 in47 sn2 21220659078919380.000000
Rwneg47_3 in47 sn3 21220659078919380.000000
Rwneg47_4 in47 sn4 21220659078919380.000000
Rwneg47_5 in47 sn5 22281692032865348.000000
Rwneg47_6 in47 sn6 22281692032865348.000000
Rwneg47_7 in47 sn7 22281692032865348.000000
Rwneg47_8 in47 sn8 21220659078919380.000000
Rwneg47_9 in47 sn9 21220659078919380.000000
Rwneg47_10 in47 sn10 22281692032865348.000000
Rwneg48_1 in48 sn1 22281692032865348.000000
Rwneg48_2 in48 sn2 21220659078919380.000000
Rwneg48_3 in48 sn3 22281692032865348.000000
Rwneg48_4 in48 sn4 22281692032865348.000000
Rwneg48_5 in48 sn5 21220659078919380.000000
Rwneg48_6 in48 sn6 22281692032865348.000000
Rwneg48_7 in48 sn7 21220659078919380.000000
Rwneg48_8 in48 sn8 22281692032865348.000000
Rwneg48_9 in48 sn9 22281692032865348.000000
Rwneg48_10 in48 sn10 22281692032865348.000000
Rwneg49_1 in49 sn1 21220659078919380.000000
Rwneg49_2 in49 sn2 22281692032865348.000000
Rwneg49_3 in49 sn3 22281692032865348.000000
Rwneg49_4 in49 sn4 22281692032865348.000000
Rwneg49_5 in49 sn5 22281692032865348.000000
Rwneg49_6 in49 sn6 21220659078919380.000000
Rwneg49_7 in49 sn7 21220659078919380.000000
Rwneg49_8 in49 sn8 21220659078919380.000000
Rwneg49_9 in49 sn9 22281692032865348.000000
Rwneg49_10 in49 sn10 22281692032865348.000000
Rwneg50_1 in50 sn1 22281692032865348.000000
Rwneg50_2 in50 sn2 21220659078919380.000000
Rwneg50_3 in50 sn3 22281692032865348.000000
Rwneg50_4 in50 sn4 21220659078919380.000000
Rwneg50_5 in50 sn5 22281692032865348.000000
Rwneg50_6 in50 sn6 22281692032865348.000000
Rwneg50_7 in50 sn7 21220659078919380.000000
Rwneg50_8 in50 sn8 21220659078919380.000000
Rwneg50_9 in50 sn9 22281692032865348.000000
Rwneg50_10 in50 sn10 21220659078919380.000000
Rwneg51_1 in51 sn1 21220659078919380.000000
Rwneg51_2 in51 sn2 22281692032865348.000000
Rwneg51_3 in51 sn3 22281692032865348.000000
Rwneg51_4 in51 sn4 21220659078919380.000000
Rwneg51_5 in51 sn5 22281692032865348.000000
Rwneg51_6 in51 sn6 21220659078919380.000000
Rwneg51_7 in51 sn7 22281692032865348.000000
Rwneg51_8 in51 sn8 21220659078919380.000000
Rwneg51_9 in51 sn9 22281692032865348.000000
Rwneg51_10 in51 sn10 22281692032865348.000000
Rwneg52_1 in52 sn1 22281692032865348.000000
Rwneg52_2 in52 sn2 22281692032865348.000000
Rwneg52_3 in52 sn3 21220659078919380.000000
Rwneg52_4 in52 sn4 21220659078919380.000000
Rwneg52_5 in52 sn5 22281692032865348.000000
Rwneg52_6 in52 sn6 21220659078919380.000000
Rwneg52_7 in52 sn7 22281692032865348.000000
Rwneg52_8 in52 sn8 21220659078919380.000000
Rwneg52_9 in52 sn9 22281692032865348.000000
Rwneg52_10 in52 sn10 22281692032865348.000000
Rwneg53_1 in53 sn1 22281692032865348.000000
Rwneg53_2 in53 sn2 21220659078919380.000000
Rwneg53_3 in53 sn3 22281692032865348.000000
Rwneg53_4 in53 sn4 22281692032865348.000000
Rwneg53_5 in53 sn5 21220659078919380.000000
Rwneg53_6 in53 sn6 21220659078919380.000000
Rwneg53_7 in53 sn7 22281692032865348.000000
Rwneg53_8 in53 sn8 21220659078919380.000000
Rwneg53_9 in53 sn9 22281692032865348.000000
Rwneg53_10 in53 sn10 21220659078919380.000000
Rwneg54_1 in54 sn1 22281692032865348.000000
Rwneg54_2 in54 sn2 21220659078919380.000000
Rwneg54_3 in54 sn3 21220659078919380.000000
Rwneg54_4 in54 sn4 21220659078919380.000000
Rwneg54_5 in54 sn5 22281692032865348.000000
Rwneg54_6 in54 sn6 21220659078919380.000000
Rwneg54_7 in54 sn7 22281692032865348.000000
Rwneg54_8 in54 sn8 21220659078919380.000000
Rwneg54_9 in54 sn9 22281692032865348.000000
Rwneg54_10 in54 sn10 22281692032865348.000000
Rwneg55_1 in55 sn1 21220659078919380.000000
Rwneg55_2 in55 sn2 22281692032865348.000000
Rwneg55_3 in55 sn3 22281692032865348.000000
Rwneg55_4 in55 sn4 22281692032865348.000000
Rwneg55_5 in55 sn5 22281692032865348.000000
Rwneg55_6 in55 sn6 21220659078919380.000000
Rwneg55_7 in55 sn7 21220659078919380.000000
Rwneg55_8 in55 sn8 22281692032865348.000000
Rwneg55_9 in55 sn9 21220659078919380.000000
Rwneg55_10 in55 sn10 21220659078919380.000000
Rwneg56_1 in56 sn1 22281692032865348.000000
Rwneg56_2 in56 sn2 21220659078919380.000000
Rwneg56_3 in56 sn3 21220659078919380.000000
Rwneg56_4 in56 sn4 21220659078919380.000000
Rwneg56_5 in56 sn5 21220659078919380.000000
Rwneg56_6 in56 sn6 21220659078919380.000000
Rwneg56_7 in56 sn7 22281692032865348.000000
Rwneg56_8 in56 sn8 21220659078919380.000000
Rwneg56_9 in56 sn9 22281692032865348.000000
Rwneg56_10 in56 sn10 22281692032865348.000000
Rwneg57_1 in57 sn1 22281692032865348.000000
Rwneg57_2 in57 sn2 21220659078919380.000000
Rwneg57_3 in57 sn3 21220659078919380.000000
Rwneg57_4 in57 sn4 22281692032865348.000000
Rwneg57_5 in57 sn5 22281692032865348.000000
Rwneg57_6 in57 sn6 21220659078919380.000000
Rwneg57_7 in57 sn7 22281692032865348.000000
Rwneg57_8 in57 sn8 22281692032865348.000000
Rwneg57_9 in57 sn9 21220659078919380.000000
Rwneg57_10 in57 sn10 21220659078919380.000000
Rwneg58_1 in58 sn1 22281692032865348.000000
Rwneg58_2 in58 sn2 22281692032865348.000000
Rwneg58_3 in58 sn3 21220659078919380.000000
Rwneg58_4 in58 sn4 22281692032865348.000000
Rwneg58_5 in58 sn5 21220659078919380.000000
Rwneg58_6 in58 sn6 22281692032865348.000000
Rwneg58_7 in58 sn7 21220659078919380.000000
Rwneg58_8 in58 sn8 22281692032865348.000000
Rwneg58_9 in58 sn9 22281692032865348.000000
Rwneg58_10 in58 sn10 21220659078919380.000000
Rwneg59_1 in59 sn1 22281692032865348.000000
Rwneg59_2 in59 sn2 21220659078919380.000000
Rwneg59_3 in59 sn3 21220659078919380.000000
Rwneg59_4 in59 sn4 22281692032865348.000000
Rwneg59_5 in59 sn5 21220659078919380.000000
Rwneg59_6 in59 sn6 21220659078919380.000000
Rwneg59_7 in59 sn7 22281692032865348.000000
Rwneg59_8 in59 sn8 21220659078919380.000000
Rwneg59_9 in59 sn9 22281692032865348.000000
Rwneg59_10 in59 sn10 21220659078919380.000000
Rwneg60_1 in60 sn1 21220659078919380.000000
Rwneg60_2 in60 sn2 21220659078919380.000000
Rwneg60_3 in60 sn3 21220659078919380.000000
Rwneg60_4 in60 sn4 22281692032865348.000000
Rwneg60_5 in60 sn5 22281692032865348.000000
Rwneg60_6 in60 sn6 22281692032865348.000000
Rwneg60_7 in60 sn7 21220659078919380.000000
Rwneg60_8 in60 sn8 22281692032865348.000000
Rwneg60_9 in60 sn9 21220659078919380.000000
Rwneg60_10 in60 sn10 21220659078919380.000000
Rwneg61_1 in61 sn1 21220659078919380.000000
Rwneg61_2 in61 sn2 21220659078919380.000000
Rwneg61_3 in61 sn3 22281692032865348.000000
Rwneg61_4 in61 sn4 22281692032865348.000000
Rwneg61_5 in61 sn5 21220659078919380.000000
Rwneg61_6 in61 sn6 21220659078919380.000000
Rwneg61_7 in61 sn7 22281692032865348.000000
Rwneg61_8 in61 sn8 21220659078919380.000000
Rwneg61_9 in61 sn9 21220659078919380.000000
Rwneg61_10 in61 sn10 22281692032865348.000000
Rwneg62_1 in62 sn1 22281692032865348.000000
Rwneg62_2 in62 sn2 21220659078919380.000000
Rwneg62_3 in62 sn3 21220659078919380.000000
Rwneg62_4 in62 sn4 22281692032865348.000000
Rwneg62_5 in62 sn5 22281692032865348.000000
Rwneg62_6 in62 sn6 22281692032865348.000000
Rwneg62_7 in62 sn7 21220659078919380.000000
Rwneg62_8 in62 sn8 21220659078919380.000000
Rwneg62_9 in62 sn9 21220659078919380.000000
Rwneg62_10 in62 sn10 22281692032865348.000000
Rwneg63_1 in63 sn1 21220659078919380.000000
Rwneg63_2 in63 sn2 21220659078919380.000000
Rwneg63_3 in63 sn3 22281692032865348.000000
Rwneg63_4 in63 sn4 22281692032865348.000000
Rwneg63_5 in63 sn5 22281692032865348.000000
Rwneg63_6 in63 sn6 21220659078919380.000000
Rwneg63_7 in63 sn7 21220659078919380.000000
Rwneg63_8 in63 sn8 21220659078919380.000000
Rwneg63_9 in63 sn9 22281692032865348.000000
Rwneg63_10 in63 sn10 22281692032865348.000000
Rwneg64_1 in64 sn1 22281692032865348.000000
Rwneg64_2 in64 sn2 22281692032865348.000000
Rwneg64_3 in64 sn3 22281692032865348.000000
Rwneg64_4 in64 sn4 22281692032865348.000000
Rwneg64_5 in64 sn5 21220659078919380.000000
Rwneg64_6 in64 sn6 22281692032865348.000000
Rwneg64_7 in64 sn7 22281692032865348.000000
Rwneg64_8 in64 sn8 22281692032865348.000000
Rwneg64_9 in64 sn9 22281692032865348.000000
Rwneg64_10 in64 sn10 22281692032865348.000000
Rwneg65_1 in65 sn1 21220659078919380.000000
Rwneg65_2 in65 sn2 22281692032865348.000000
Rwneg65_3 in65 sn3 21220659078919380.000000
Rwneg65_4 in65 sn4 22281692032865348.000000
Rwneg65_5 in65 sn5 22281692032865348.000000
Rwneg65_6 in65 sn6 22281692032865348.000000
Rwneg65_7 in65 sn7 22281692032865348.000000
Rwneg65_8 in65 sn8 21220659078919380.000000
Rwneg65_9 in65 sn9 21220659078919380.000000
Rwneg65_10 in65 sn10 22281692032865348.000000
Rwneg66_1 in66 sn1 22281692032865348.000000
Rwneg66_2 in66 sn2 21220659078919380.000000
Rwneg66_3 in66 sn3 22281692032865348.000000
Rwneg66_4 in66 sn4 21220659078919380.000000
Rwneg66_5 in66 sn5 21220659078919380.000000
Rwneg66_6 in66 sn6 22281692032865348.000000
Rwneg66_7 in66 sn7 21220659078919380.000000
Rwneg66_8 in66 sn8 21220659078919380.000000
Rwneg66_9 in66 sn9 22281692032865348.000000
Rwneg66_10 in66 sn10 22281692032865348.000000
Rwneg67_1 in67 sn1 22281692032865348.000000
Rwneg67_2 in67 sn2 21220659078919380.000000
Rwneg67_3 in67 sn3 21220659078919380.000000
Rwneg67_4 in67 sn4 22281692032865348.000000
Rwneg67_5 in67 sn5 22281692032865348.000000
Rwneg67_6 in67 sn6 21220659078919380.000000
Rwneg67_7 in67 sn7 21220659078919380.000000
Rwneg67_8 in67 sn8 22281692032865348.000000
Rwneg67_9 in67 sn9 22281692032865348.000000
Rwneg67_10 in67 sn10 22281692032865348.000000
Rwneg68_1 in68 sn1 21220659078919380.000000
Rwneg68_2 in68 sn2 21220659078919380.000000
Rwneg68_3 in68 sn3 21220659078919380.000000
Rwneg68_4 in68 sn4 22281692032865348.000000
Rwneg68_5 in68 sn5 22281692032865348.000000
Rwneg68_6 in68 sn6 21220659078919380.000000
Rwneg68_7 in68 sn7 22281692032865348.000000
Rwneg68_8 in68 sn8 21220659078919380.000000
Rwneg68_9 in68 sn9 22281692032865348.000000
Rwneg68_10 in68 sn10 22281692032865348.000000
Rwneg69_1 in69 sn1 22281692032865348.000000
Rwneg69_2 in69 sn2 21220659078919380.000000
Rwneg69_3 in69 sn3 22281692032865348.000000
Rwneg69_4 in69 sn4 21220659078919380.000000
Rwneg69_5 in69 sn5 22281692032865348.000000
Rwneg69_6 in69 sn6 21220659078919380.000000
Rwneg69_7 in69 sn7 21220659078919380.000000
Rwneg69_8 in69 sn8 22281692032865348.000000
Rwneg69_9 in69 sn9 21220659078919380.000000
Rwneg69_10 in69 sn10 21220659078919380.000000
Rwneg70_1 in70 sn1 22281692032865348.000000
Rwneg70_2 in70 sn2 21220659078919380.000000
Rwneg70_3 in70 sn3 21220659078919380.000000
Rwneg70_4 in70 sn4 22281692032865348.000000
Rwneg70_5 in70 sn5 21220659078919380.000000
Rwneg70_6 in70 sn6 22281692032865348.000000
Rwneg70_7 in70 sn7 21220659078919380.000000
Rwneg70_8 in70 sn8 21220659078919380.000000
Rwneg70_9 in70 sn9 22281692032865348.000000
Rwneg70_10 in70 sn10 21220659078919380.000000
Rwneg71_1 in71 sn1 22281692032865348.000000
Rwneg71_2 in71 sn2 21220659078919380.000000
Rwneg71_3 in71 sn3 21220659078919380.000000
Rwneg71_4 in71 sn4 21220659078919380.000000
Rwneg71_5 in71 sn5 22281692032865348.000000
Rwneg71_6 in71 sn6 21220659078919380.000000
Rwneg71_7 in71 sn7 22281692032865348.000000
Rwneg71_8 in71 sn8 22281692032865348.000000
Rwneg71_9 in71 sn9 21220659078919380.000000
Rwneg71_10 in71 sn10 21220659078919380.000000
Rwneg72_1 in72 sn1 22281692032865348.000000
Rwneg72_2 in72 sn2 21220659078919380.000000
Rwneg72_3 in72 sn3 21220659078919380.000000
Rwneg72_4 in72 sn4 21220659078919380.000000
Rwneg72_5 in72 sn5 21220659078919380.000000
Rwneg72_6 in72 sn6 22281692032865348.000000
Rwneg72_7 in72 sn7 22281692032865348.000000
Rwneg72_8 in72 sn8 21220659078919380.000000
Rwneg72_9 in72 sn9 22281692032865348.000000
Rwneg72_10 in72 sn10 22281692032865348.000000
Rwneg73_1 in73 sn1 21220659078919380.000000
Rwneg73_2 in73 sn2 21220659078919380.000000
Rwneg73_3 in73 sn3 22281692032865348.000000
Rwneg73_4 in73 sn4 21220659078919380.000000
Rwneg73_5 in73 sn5 21220659078919380.000000
Rwneg73_6 in73 sn6 22281692032865348.000000
Rwneg73_7 in73 sn7 22281692032865348.000000
Rwneg73_8 in73 sn8 22281692032865348.000000
Rwneg73_9 in73 sn9 21220659078919380.000000
Rwneg73_10 in73 sn10 21220659078919380.000000
Rwneg74_1 in74 sn1 22281692032865348.000000
Rwneg74_2 in74 sn2 22281692032865348.000000
Rwneg74_3 in74 sn3 22281692032865348.000000
Rwneg74_4 in74 sn4 21220659078919380.000000
Rwneg74_5 in74 sn5 21220659078919380.000000
Rwneg74_6 in74 sn6 21220659078919380.000000
Rwneg74_7 in74 sn7 21220659078919380.000000
Rwneg74_8 in74 sn8 22281692032865348.000000
Rwneg74_9 in74 sn9 21220659078919380.000000
Rwneg74_10 in74 sn10 22281692032865348.000000
Rwneg75_1 in75 sn1 22281692032865348.000000
Rwneg75_2 in75 sn2 22281692032865348.000000
Rwneg75_3 in75 sn3 22281692032865348.000000
Rwneg75_4 in75 sn4 21220659078919380.000000
Rwneg75_5 in75 sn5 21220659078919380.000000
Rwneg75_6 in75 sn6 22281692032865348.000000
Rwneg75_7 in75 sn7 22281692032865348.000000
Rwneg75_8 in75 sn8 21220659078919380.000000
Rwneg75_9 in75 sn9 22281692032865348.000000
Rwneg75_10 in75 sn10 21220659078919380.000000
Rwneg76_1 in76 sn1 22281692032865348.000000
Rwneg76_2 in76 sn2 21220659078919380.000000
Rwneg76_3 in76 sn3 21220659078919380.000000
Rwneg76_4 in76 sn4 21220659078919380.000000
Rwneg76_5 in76 sn5 21220659078919380.000000
Rwneg76_6 in76 sn6 22281692032865348.000000
Rwneg76_7 in76 sn7 22281692032865348.000000
Rwneg76_8 in76 sn8 22281692032865348.000000
Rwneg76_9 in76 sn9 22281692032865348.000000
Rwneg76_10 in76 sn10 21220659078919380.000000
Rwneg77_1 in77 sn1 22281692032865348.000000
Rwneg77_2 in77 sn2 22281692032865348.000000
Rwneg77_3 in77 sn3 21220659078919380.000000
Rwneg77_4 in77 sn4 22281692032865348.000000
Rwneg77_5 in77 sn5 21220659078919380.000000
Rwneg77_6 in77 sn6 21220659078919380.000000
Rwneg77_7 in77 sn7 21220659078919380.000000
Rwneg77_8 in77 sn8 22281692032865348.000000
Rwneg77_9 in77 sn9 22281692032865348.000000
Rwneg77_10 in77 sn10 22281692032865348.000000
Rwneg78_1 in78 sn1 21220659078919380.000000
Rwneg78_2 in78 sn2 22281692032865348.000000
Rwneg78_3 in78 sn3 21220659078919380.000000
Rwneg78_4 in78 sn4 21220659078919380.000000
Rwneg78_5 in78 sn5 22281692032865348.000000
Rwneg78_6 in78 sn6 21220659078919380.000000
Rwneg78_7 in78 sn7 22281692032865348.000000
Rwneg78_8 in78 sn8 22281692032865348.000000
Rwneg78_9 in78 sn9 22281692032865348.000000
Rwneg78_10 in78 sn10 21220659078919380.000000
Rwneg79_1 in79 sn1 22281692032865348.000000
Rwneg79_2 in79 sn2 21220659078919380.000000
Rwneg79_3 in79 sn3 21220659078919380.000000
Rwneg79_4 in79 sn4 22281692032865348.000000
Rwneg79_5 in79 sn5 21220659078919380.000000
Rwneg79_6 in79 sn6 21220659078919380.000000
Rwneg79_7 in79 sn7 22281692032865348.000000
Rwneg79_8 in79 sn8 21220659078919380.000000
Rwneg79_9 in79 sn9 22281692032865348.000000
Rwneg79_10 in79 sn10 22281692032865348.000000
Rwneg80_1 in80 sn1 22281692032865348.000000
Rwneg80_2 in80 sn2 21220659078919380.000000
Rwneg80_3 in80 sn3 22281692032865348.000000
Rwneg80_4 in80 sn4 21220659078919380.000000
Rwneg80_5 in80 sn5 22281692032865348.000000
Rwneg80_6 in80 sn6 21220659078919380.000000
Rwneg80_7 in80 sn7 21220659078919380.000000
Rwneg80_8 in80 sn8 22281692032865348.000000
Rwneg80_9 in80 sn9 21220659078919380.000000
Rwneg80_10 in80 sn10 22281692032865348.000000
Rwneg81_1 in81 sn1 21220659078919380.000000
Rwneg81_2 in81 sn2 21220659078919380.000000
Rwneg81_3 in81 sn3 22281692032865348.000000
Rwneg81_4 in81 sn4 21220659078919380.000000
Rwneg81_5 in81 sn5 21220659078919380.000000
Rwneg81_6 in81 sn6 22281692032865348.000000
Rwneg81_7 in81 sn7 21220659078919380.000000
Rwneg81_8 in81 sn8 21220659078919380.000000
Rwneg81_9 in81 sn9 22281692032865348.000000
Rwneg81_10 in81 sn10 22281692032865348.000000
Rwneg82_1 in82 sn1 21220659078919380.000000
Rwneg82_2 in82 sn2 21220659078919380.000000
Rwneg82_3 in82 sn3 21220659078919380.000000
Rwneg82_4 in82 sn4 21220659078919380.000000
Rwneg82_5 in82 sn5 22281692032865348.000000
Rwneg82_6 in82 sn6 22281692032865348.000000
Rwneg82_7 in82 sn7 21220659078919380.000000
Rwneg82_8 in82 sn8 22281692032865348.000000
Rwneg82_9 in82 sn9 22281692032865348.000000
Rwneg82_10 in82 sn10 21220659078919380.000000
Rwneg83_1 in83 sn1 22281692032865348.000000
Rwneg83_2 in83 sn2 21220659078919380.000000
Rwneg83_3 in83 sn3 21220659078919380.000000
Rwneg83_4 in83 sn4 22281692032865348.000000
Rwneg83_5 in83 sn5 22281692032865348.000000
Rwneg83_6 in83 sn6 22281692032865348.000000
Rwneg83_7 in83 sn7 21220659078919380.000000
Rwneg83_8 in83 sn8 22281692032865348.000000
Rwneg83_9 in83 sn9 22281692032865348.000000
Rwneg83_10 in83 sn10 22281692032865348.000000
Rwneg84_1 in84 sn1 21220659078919380.000000
Rwneg84_2 in84 sn2 22281692032865348.000000
Rwneg84_3 in84 sn3 22281692032865348.000000
Rwneg84_4 in84 sn4 22281692032865348.000000
Rwneg84_5 in84 sn5 21220659078919380.000000
Rwneg84_6 in84 sn6 22281692032865348.000000
Rwneg84_7 in84 sn7 22281692032865348.000000
Rwneg84_8 in84 sn8 21220659078919380.000000
Rwneg84_9 in84 sn9 22281692032865348.000000
Rwneg84_10 in84 sn10 21220659078919380.000000
Rwneg85_1 in85 sn1 21220659078919380.000000
Rwneg85_2 in85 sn2 21220659078919380.000000
Rwneg85_3 in85 sn3 21220659078919380.000000
Rwneg85_4 in85 sn4 22281692032865348.000000
Rwneg85_5 in85 sn5 22281692032865348.000000
Rwneg85_6 in85 sn6 22281692032865348.000000
Rwneg85_7 in85 sn7 21220659078919380.000000
Rwneg85_8 in85 sn8 22281692032865348.000000
Rwneg85_9 in85 sn9 22281692032865348.000000
Rwneg85_10 in85 sn10 21220659078919380.000000
Rwneg86_1 in86 sn1 21220659078919380.000000
Rwneg86_2 in86 sn2 21220659078919380.000000
Rwneg86_3 in86 sn3 22281692032865348.000000
Rwneg86_4 in86 sn4 22281692032865348.000000
Rwneg86_5 in86 sn5 21220659078919380.000000
Rwneg86_6 in86 sn6 22281692032865348.000000
Rwneg86_7 in86 sn7 22281692032865348.000000
Rwneg86_8 in86 sn8 22281692032865348.000000
Rwneg86_9 in86 sn9 21220659078919380.000000
Rwneg86_10 in86 sn10 22281692032865348.000000
Rwneg87_1 in87 sn1 22281692032865348.000000
Rwneg87_2 in87 sn2 21220659078919380.000000
Rwneg87_3 in87 sn3 22281692032865348.000000
Rwneg87_4 in87 sn4 22281692032865348.000000
Rwneg87_5 in87 sn5 22281692032865348.000000
Rwneg87_6 in87 sn6 21220659078919380.000000
Rwneg87_7 in87 sn7 22281692032865348.000000
Rwneg87_8 in87 sn8 21220659078919380.000000
Rwneg87_9 in87 sn9 22281692032865348.000000
Rwneg87_10 in87 sn10 21220659078919380.000000
Rwneg88_1 in88 sn1 22281692032865348.000000
Rwneg88_2 in88 sn2 22281692032865348.000000
Rwneg88_3 in88 sn3 21220659078919380.000000
Rwneg88_4 in88 sn4 22281692032865348.000000
Rwneg88_5 in88 sn5 21220659078919380.000000
Rwneg88_6 in88 sn6 21220659078919380.000000
Rwneg88_7 in88 sn7 22281692032865348.000000
Rwneg88_8 in88 sn8 21220659078919380.000000
Rwneg88_9 in88 sn9 22281692032865348.000000
Rwneg88_10 in88 sn10 21220659078919380.000000
Rwneg89_1 in89 sn1 21220659078919380.000000
Rwneg89_2 in89 sn2 22281692032865348.000000
Rwneg89_3 in89 sn3 21220659078919380.000000
Rwneg89_4 in89 sn4 21220659078919380.000000
Rwneg89_5 in89 sn5 22281692032865348.000000
Rwneg89_6 in89 sn6 22281692032865348.000000
Rwneg89_7 in89 sn7 22281692032865348.000000
Rwneg89_8 in89 sn8 21220659078919380.000000
Rwneg89_9 in89 sn9 21220659078919380.000000
Rwneg89_10 in89 sn10 21220659078919380.000000
Rwneg90_1 in90 sn1 22281692032865348.000000
Rwneg90_2 in90 sn2 21220659078919380.000000
Rwneg90_3 in90 sn3 22281692032865348.000000
Rwneg90_4 in90 sn4 21220659078919380.000000
Rwneg90_5 in90 sn5 22281692032865348.000000
Rwneg90_6 in90 sn6 21220659078919380.000000
Rwneg90_7 in90 sn7 22281692032865348.000000
Rwneg90_8 in90 sn8 22281692032865348.000000
Rwneg90_9 in90 sn9 22281692032865348.000000
Rwneg90_10 in90 sn10 21220659078919380.000000
Rwneg91_1 in91 sn1 22281692032865348.000000
Rwneg91_2 in91 sn2 22281692032865348.000000
Rwneg91_3 in91 sn3 21220659078919380.000000
Rwneg91_4 in91 sn4 22281692032865348.000000
Rwneg91_5 in91 sn5 22281692032865348.000000
Rwneg91_6 in91 sn6 22281692032865348.000000
Rwneg91_7 in91 sn7 21220659078919380.000000
Rwneg91_8 in91 sn8 21220659078919380.000000
Rwneg91_9 in91 sn9 22281692032865348.000000
Rwneg91_10 in91 sn10 21220659078919380.000000
Rwneg92_1 in92 sn1 22281692032865348.000000
Rwneg92_2 in92 sn2 22281692032865348.000000
Rwneg92_3 in92 sn3 22281692032865348.000000
Rwneg92_4 in92 sn4 22281692032865348.000000
Rwneg92_5 in92 sn5 22281692032865348.000000
Rwneg92_6 in92 sn6 22281692032865348.000000
Rwneg92_7 in92 sn7 21220659078919380.000000
Rwneg92_8 in92 sn8 22281692032865348.000000
Rwneg92_9 in92 sn9 22281692032865348.000000
Rwneg92_10 in92 sn10 22281692032865348.000000
Rwneg93_1 in93 sn1 22281692032865348.000000
Rwneg93_2 in93 sn2 21220659078919380.000000
Rwneg93_3 in93 sn3 22281692032865348.000000
Rwneg93_4 in93 sn4 22281692032865348.000000
Rwneg93_5 in93 sn5 22281692032865348.000000
Rwneg93_6 in93 sn6 21220659078919380.000000
Rwneg93_7 in93 sn7 21220659078919380.000000
Rwneg93_8 in93 sn8 21220659078919380.000000
Rwneg93_9 in93 sn9 22281692032865348.000000
Rwneg93_10 in93 sn10 21220659078919380.000000
Rwneg94_1 in94 sn1 21220659078919380.000000
Rwneg94_2 in94 sn2 22281692032865348.000000
Rwneg94_3 in94 sn3 22281692032865348.000000
Rwneg94_4 in94 sn4 22281692032865348.000000
Rwneg94_5 in94 sn5 21220659078919380.000000
Rwneg94_6 in94 sn6 21220659078919380.000000
Rwneg94_7 in94 sn7 22281692032865348.000000
Rwneg94_8 in94 sn8 22281692032865348.000000
Rwneg94_9 in94 sn9 22281692032865348.000000
Rwneg94_10 in94 sn10 21220659078919380.000000
Rwneg95_1 in95 sn1 21220659078919380.000000
Rwneg95_2 in95 sn2 22281692032865348.000000
Rwneg95_3 in95 sn3 21220659078919380.000000
Rwneg95_4 in95 sn4 22281692032865348.000000
Rwneg95_5 in95 sn5 22281692032865348.000000
Rwneg95_6 in95 sn6 21220659078919380.000000
Rwneg95_7 in95 sn7 22281692032865348.000000
Rwneg95_8 in95 sn8 22281692032865348.000000
Rwneg95_9 in95 sn9 21220659078919380.000000
Rwneg95_10 in95 sn10 21220659078919380.000000
Rwneg96_1 in96 sn1 21220659078919380.000000
Rwneg96_2 in96 sn2 22281692032865348.000000
Rwneg96_3 in96 sn3 21220659078919380.000000
Rwneg96_4 in96 sn4 22281692032865348.000000
Rwneg96_5 in96 sn5 21220659078919380.000000
Rwneg96_6 in96 sn6 22281692032865348.000000
Rwneg96_7 in96 sn7 21220659078919380.000000
Rwneg96_8 in96 sn8 22281692032865348.000000
Rwneg96_9 in96 sn9 21220659078919380.000000
Rwneg96_10 in96 sn10 22281692032865348.000000
Rwneg97_1 in97 sn1 22281692032865348.000000
Rwneg97_2 in97 sn2 21220659078919380.000000
Rwneg97_3 in97 sn3 21220659078919380.000000
Rwneg97_4 in97 sn4 22281692032865348.000000
Rwneg97_5 in97 sn5 21220659078919380.000000
Rwneg97_6 in97 sn6 21220659078919380.000000
Rwneg97_7 in97 sn7 22281692032865348.000000
Rwneg97_8 in97 sn8 21220659078919380.000000
Rwneg97_9 in97 sn9 21220659078919380.000000
Rwneg97_10 in97 sn10 21220659078919380.000000
Rwneg98_1 in98 sn1 21220659078919380.000000
Rwneg98_2 in98 sn2 22281692032865348.000000
Rwneg98_3 in98 sn3 22281692032865348.000000
Rwneg98_4 in98 sn4 22281692032865348.000000
Rwneg98_5 in98 sn5 21220659078919380.000000
Rwneg98_6 in98 sn6 21220659078919380.000000
Rwneg98_7 in98 sn7 21220659078919380.000000
Rwneg98_8 in98 sn8 21220659078919380.000000
Rwneg98_9 in98 sn9 21220659078919380.000000
Rwneg98_10 in98 sn10 22281692032865348.000000
Rwneg99_1 in99 sn1 21220659078919380.000000
Rwneg99_2 in99 sn2 21220659078919380.000000
Rwneg99_3 in99 sn3 21220659078919380.000000
Rwneg99_4 in99 sn4 22281692032865348.000000
Rwneg99_5 in99 sn5 21220659078919380.000000
Rwneg99_6 in99 sn6 21220659078919380.000000
Rwneg99_7 in99 sn7 21220659078919380.000000
Rwneg99_8 in99 sn8 21220659078919380.000000
Rwneg99_9 in99 sn9 22281692032865348.000000
Rwneg99_10 in99 sn10 22281692032865348.000000
Rwneg100_1 in100 sn1 22281692032865348.000000
Rwneg100_2 in100 sn2 22281692032865348.000000
Rwneg100_3 in100 sn3 21220659078919380.000000
Rwneg100_4 in100 sn4 21220659078919380.000000
Rwneg100_5 in100 sn5 22281692032865348.000000
Rwneg100_6 in100 sn6 21220659078919380.000000
Rwneg100_7 in100 sn7 22281692032865348.000000
Rwneg100_8 in100 sn8 21220659078919380.000000
Rwneg100_9 in100 sn9 21220659078919380.000000
Rwneg100_10 in100 sn10 22281692032865348.000000


**********Positive Biases****************

Rbpos1 vdd sp1 21220659078919380.000000
Rbpos2 vdd sp2 21220659078919380.000000
Rbpos3 vdd sp3 21220659078919380.000000
Rbpos4 vdd sp4 21220659078919380.000000
Rbpos5 vdd sp5 21220659078919380.000000
Rbpos6 vdd sp6 21220659078919380.000000
Rbpos7 vdd sp7 21220659078919380.000000
Rbpos8 vdd sp8 21220659078919380.000000
Rbpos9 vdd sp9 21220659078919380.000000
Rbpos10 vdd sp10 21220659078919380.000000


**********Negative Biases****************

Rbneg1 vss sn1 22281692032865348.000000
Rbneg2 vss sn2 22281692032865348.000000
Rbneg3 vss sn3 22281692032865348.000000
Rbneg4 vss sn4 22281692032865348.000000
Rbneg5 vss sn5 22281692032865348.000000
Rbneg6 vss sn6 22281692032865348.000000
Rbneg7 vss sn7 22281692032865348.000000
Rbneg8 vss sn8 22281692032865348.000000
Rbneg9 vss sn9 22281692032865348.000000
Rbneg10 vss sn10 22281692032865348.000000


**********Weight Differntial Op-AMPS****************

XDIFFw1 sp1 sn1 xin1 diff2
XDIFFw2 sp2 sn2 xin2 diff2
XDIFFw3 sp3 sn3 xin3 diff2
XDIFFw4 sp4 sn4 xin4 diff2
XDIFFw5 sp5 sn5 xin5 diff2
XDIFFw6 sp6 sn6 xin6 diff2
XDIFFw7 sp7 sn7 xin7 diff2
XDIFFw8 sp8 sn8 xin8 diff2
XDIFFw9 sp9 sn9 xin9 diff2
XDIFFw10 sp10 sn10 xin10 diff2


**********neurons****************

Xsig1 xin1 out1 vdd 0 neuron
Xsig2 xin2 out2 vdd 0 neuron
Xsig3 xin3 out3 vdd 0 neuron
Xsig4 xin4 out4 vdd 0 neuron
Xsig5 xin5 out5 vdd 0 neuron
Xsig6 xin6 out6 vdd 0 neuron
Xsig7 xin7 out7 vdd 0 neuron
Xsig8 xin8 out8 vdd 0 neuron
Xsig9 xin9 out9 vdd 0 neuron
Xsig10 xin10 out10 vdd 0 neuron
.ENDS layer2